.subckt data_reg_bank clk rst x_in_0 x_in_1 x_in_2 x_in_3 y_in_0 y_in_1 y_in_2 y_in_3 x_out_0 x_out_1 x_out_2 x_out_3 x_out_b_0 x_out_b_1 x_out_b_2 x_out_b_3 y_out_0 y_out_1 y_out_2 y_out_3 y_out_b_0 y_out_b_1 y_out_b_2 y_out_b_3 clk_div4_out clk_div4_out_b vdd vss


** Library name: final_project_local
** Cell name: data_reg_bank
** View name: av_extracted
c1 vdd vss 181.257e-18
c2 clk vss 101.165e-18
c3 rst vss 256.643e-18
c4 x_in_0 vss 9.56674e-18
c5 x_in_1 vss 8.92083e-18
c6 x_in_2 vss 9.56674e-18
c7 x_in_3 vss 8.94641e-18
c8 y_in_0 vss 438.192e-18
c9 y_in_1 vss 494.358e-18
c10 y_in_2 vss 494.369e-18
c11 y_in_3 vss 438.452e-18
c12 clk_div4_out vss 121.735e-18
c13 clk_div4_out_b vss 157.065e-18
c14 x_out_0 vss 187.294e-18
c15 x_out_1 vss 186.127e-18
c16 x_out_2 vss 187.616e-18
c17 x_out_3 vss 185.948e-18
c18 x_out_b_0 vss 155.079e-18
c19 x_out_b_1 vss 155.078e-18
c20 x_out_b_2 vss 155.079e-18
c21 x_out_b_3 vss 155.079e-18
c22 y_out_0 vss 35.8556e-18
c23 y_out_1 vss 38.8088e-18
c24 y_out_2 vss 38.807e-18
c25 y_out_3 vss 37.944e-18
c26 y_out_b_0 vss 105.536e-18
c27 y_out_b_1 vss 107.227e-18
c28 y_out_b_2 vss 107.229e-18
c29 y_out_b_3 vss 107.227e-18
c30 net7 vss 20.0926e-18
c31 net11 vss 21.793e-18
c32 net9 vss 31.6438e-18
c33 net10 vss 29.561e-18
c34 net3 vss 21.4174e-18
c35 net4 vss 16.5107e-18
c36 avs88 vss 195.269e-18
c37 i0__net10 vss 21.3377e-18
c38 i0__net9 vss 21.6046e-18
c39 i0__net8 vss 57.1298e-18
c40 i0__net11 vss 32.9291e-18
c41 i0__net1 vss 31.0739e-18
c42 i0__net7 vss 82.7703e-18
c43 i0__net6 vss 16.52e-18
c44 i0__net3 vss 28.9417e-18
c45 i0__i2__net5 vss 17.1191e-18
c46 i0__i2__net4 vss 113.401e-18
c47 i0__i2__net1 vss 18.0509e-18
c48 i0__i2__net2 vss 117.361e-18
c49 i0__i3__net5 vss 23.6687e-18
c50 i0__i3__net4 vss 109.189e-18
c51 i0__i3__net1 vss 26.5256e-18
c52 i0__i3__net2 vss 111.841e-18
c53 i7__net5 vss 19.924e-18
c54 i7__net4 vss 114.572e-18
c55 i7__net1 vss 20.8659e-18
c56 i7__net2 vss 114.023e-18
c57 i1__net5 vss 17.5366e-18
c58 i1__net4 vss 112.638e-18
c59 i1__net1 vss 18.4343e-18
c60 i1__net2 vss 115.972e-18
c61 i4__net5 vss 18.5658e-18
c62 i4__net4 vss 114.045e-18
c63 i4__net1 vss 18.8969e-18
c64 i4__net2 vss 115.452e-18
c65 i3__net5 vss 18.7278e-18
c66 i3__net4 vss 113.256e-18
c67 i3__net1 vss 19.4125e-18
c68 i3__net2 vss 116.298e-18
c69 i6__net5 vss 24.425e-18
c70 i6__net4 vss 109.694e-18
c71 i6__net1 vss 26.2872e-18
c72 i6__net2 vss 109.307e-18
c73 i2__net5 vss 24.0926e-18
c74 i2__net4 vss 108.727e-18
c75 i2__net1 vss 26.1676e-18
c76 i2__net2 vss 110.07e-18
c77 i5__net5 vss 24.4221e-18
c78 i5__net4 vss 108.151e-18
c79 i5__net1 vss 26.2874e-18
c80 i5__net2 vss 108.418e-18
c81 i8__net5 vss 24.0926e-18
c82 i8__net4 vss 108.001e-18
c83 i8__net1 vss 26.1676e-18
c84 i8__net2 vss 109.577e-18
c85 n15__net7 vss 23.915e-18
c86 n5__net11 vss 24.7755e-18
c87 n4__y_out_b_3 vss 27.6313e-18
c88 n1__y_out_b_2 vss 27.5946e-18
c89 n4__y_out_b_1 vss 27.6313e-18
c90 n1__y_out_b_0 vss 27.5633e-18
c91 n16__net7 vss 18.865e-18
c92 n17__net11 vss 19.1502e-18
c93 n18__net7 vss 18.9853e-18
c94 n19__net11 vss 18.7421e-18
c95 n6__i7__net4 vss 29.9865e-18
c96 n4__i6__net4 vss 31.4048e-18
c97 n6__i4__net4 vss 29.9865e-18
c98 n4__i5__net4 vss 31.4048e-18
c99 n20__net7 vss 19.3126e-18
c100 n21__net11 vss 19.0498e-18
c101 n22__net7 vss 18.8717e-18
c102 n23__net11 vss 18.722e-18
c103 n5__i7__net5 vss 23.0202e-18
c104 n5__i4__net5 vss 23.0202e-18
c105 n14__net7 vss 24.7145e-18
c106 n24__net11 vss 24.3573e-18
c107 n6__i7__net5 vss 26.3916e-18
c108 n7__i6__net5 vss 26.3689e-18
c109 n6__i4__net5 vss 26.3916e-18
c110 n7__i5__net5 vss 26.3689e-18
c111 n29__net4 vss 25.9388e-18
c112 n4__net11 vss 30.1198e-18
c113 n21__net4 vss 16.1491e-18
c114 n23__net4 vss 16.1491e-18
c115 n25__net4 vss 16.1491e-18
c116 n27__net4 vss 16.1491e-18
c117 n41__net4 vss 17.9049e-18
c118 n43__net4 vss 14.9656e-18
c119 n4__net7 vss 28.7891e-18
c120 n2__i7__net4 vss 30.2474e-18
c121 n3__i6__net4 vss 29.744e-18
c122 n2__i4__net4 vss 30.2523e-18
c123 n3__i5__net4 vss 29.744e-18
c124 n45__net4 vss 19.1736e-18
c125 n47__net4 vss 15.0491e-18
c126 n48__net4 vss 25.6194e-18
c127 n50__net9 vss 16.6823e-18
c128 n52__net9 vss 16.6235e-18
c129 n54__net9 vss 16.6823e-18
c130 n56__net9 vss 16.6235e-18
c131 n33__rst vss 21.4431e-18
c132 n6__i0__net11 vss 37.6501e-18
c133 n34__rst vss 19.5045e-18
c134 n5__i7__net1 vss 26.8189e-18
c135 n5__i4__net1 vss 26.819e-18
c136 n15__i0__net8 vss 40.9128e-18
c137 n36__rst vss 18.8109e-18
c138 n6__i7__net1 vss 24.793e-18
c139 n7__i6__net1 vss 24.7685e-18
c140 n6__i4__net1 vss 24.7933e-18
c141 n7__i5__net1 vss 24.7688e-18
c142 n38__rst vss 15.7863e-18
c143 n40__rst vss 17.701e-18
c144 n5__i0__net10 vss 28.0174e-18
c145 n32__rst vss 21.8197e-18
c146 n5__i0__net9 vss 29.3676e-18
c147 n4__i0__net9 vss 27.8375e-18
c148 n2__i0__net11 vss 50.4804e-18
c149 n2__i7__net2 vss 28.9261e-18
c150 n3__i6__net2 vss 28.2135e-18
c151 n2__i4__net2 vss 28.9261e-18
c152 n3__i5__net2 vss 28.2135e-18
c153 n4__i0__net10 vss 30.6142e-18
c154 n10__i0__net8 vss 28.7659e-18
c155 n42__net10 vss 17.3312e-18
c156 n44__net10 vss 17.3312e-18
c157 n46__net10 vss 17.3312e-18
c158 n48__net10 vss 17.3312e-18
c159 n17__i0__net1 vss 26.7532e-18
c160 n6__i0__net8 vss 25.161e-18
c161 n6__i0__i2__net4 vss 29.6175e-18
c162 n4__i0__i3__net4 vss 31.2159e-18
c163 n4__x_out_b_3 vss 30.4966e-18
c164 n1__x_out_b_2 vss 30.4937e-18
c165 n4__x_out_b_1 vss 30.4966e-18
c166 n1__x_out_b_0 vss 30.4937e-18
c167 n5__i0__i2__net5 vss 21.9368e-18
c168 n6__i1__net4 vss 29.531e-18
c169 n4__i2__net4 vss 30.9417e-18
c170 n6__i3__net4 vss 29.5733e-18
c171 n4__i8__net4 vss 30.9417e-18
c172 n6__i0__i2__net5 vss 26.1816e-18
c173 n7__i0__i3__net5 vss 25.5608e-18
c174 n5__i1__net5 vss 22.6899e-18
c175 n5__i3__net5 vss 22.6899e-18
c176 n3__i0__net6 vss 16.3177e-18
c177 n6__i1__net5 vss 26.4304e-18
c178 n7__i2__net5 vss 26.4079e-18
c179 n6__i3__net5 vss 26.4304e-18
c180 n7__i8__net5 vss 26.4079e-18
c181 n2__i0__i2__net4 vss 31.0656e-18
c182 n3__i0__i3__net4 vss 30.862e-18
c183 n3__net4 vss 16.5107e-18
c184 n5__net4 vss 16.5107e-18
c185 n7__net4 vss 16.5107e-18
c186 n2__i1__net4 vss 31.2817e-18
c187 n3__i2__net4 vss 32.2929e-18
c188 n2__i3__net4 vss 32.329e-18
c189 n3__i8__net4 vss 32.2929e-18
c190 n4__i0__net3 vss 19.1438e-18
c191 n4__i0__net1 vss 19.0215e-18
c192 n5__i0__i2__net1 vss 26.671e-18
c193 n10__net9 vss 16.953e-18
c194 n12__net9 vss 16.8941e-18
c195 n14__net9 vss 16.953e-18
c196 n16__net9 vss 16.8941e-18
c197 n6__i0__i2__net1 vss 25.2364e-18
c198 n7__i0__i3__net1 vss 25.019e-18
c199 n5__i1__net1 vss 26.2939e-18
c200 n5__i3__net1 vss 26.2939e-18
c201 n6__i1__net1 vss 25.5452e-18
c202 n7__i2__net1 vss 25.5479e-18
c203 n6__i3__net1 vss 25.5725e-18
c204 n7__i8__net1 vss 25.5479e-18
c205 n2__i0__i2__net2 vss 29.964e-18
c206 n3__i0__i3__net2 vss 28.3945e-18
c207 n2__i1__net2 vss 31.2049e-18
c208 n3__i2__net2 vss 30.5513e-18
c209 n2__i3__net2 vss 31.2468e-18
c210 n3__i8__net2 vss 30.5094e-18
c211 n5__clk vss 16.938e-18
c212 n2__i0__net7 vss 19.2894e-18
c213 n3__clk vss 20.0697e-18
c214 n1__rst vss 39.0336e-18
c215 n2__net10 vss 17.4906e-18
c216 n4__net10 vss 17.3679e-18
c217 n6__net10 vss 17.4906e-18
c218 n8__net10 vss 17.3679e-18
c219 n5__net7 vss 16.895e-18
c220 n15__net11 vss 18.0538e-18
c221 n1__y_out_b_3 vss 21.1215e-18
c222 n4__y_out_b_2 vss 21.7364e-18
c223 n1__y_out_b_1 vss 21.8171e-18
c224 n4__y_out_b_0 vss 19.3005e-18
c225 n17__net7 vss 12.4378e-18
c226 n16__net11 vss 13.7909e-18
c227 n19__net7 vss 11.8577e-18
c228 n18__net11 vss 12.7931e-18
c229 n4__i7__net4 vss 26.0708e-18
c230 n6__i6__net4 vss 23.4387e-18
c231 n4__i4__net4 vss 25.0237e-18
c232 n6__i5__net4 vss 20.7763e-18
c233 n21__net7 vss 11.8327e-18
c234 n20__net11 vss 12.6114e-18
c235 n23__net7 vss 11.8165e-18
c236 n22__net11 vss 11.9394e-18
c237 n5__i6__net5 vss 17.1572e-18
c238 n5__i5__net5 vss 15.2713e-18
c239 n24__net7 vss 16.9975e-18
c240 n14__net11 vss 19.334e-18
c241 n7__i7__net5 vss 20.2153e-18
c242 n6__i6__net5 vss 22.5411e-18
c243 n7__i4__net5 vss 22.515e-18
c244 n6__i5__net5 vss 19.3045e-18
c245 n39__net4 vss 15.914e-18
c246 n40__net4 vss 14.7545e-18
c247 n3__i7__net4 vss 68.1767e-18
c248 n2__i6__net4 vss 71.8362e-18
c249 n3__i4__net4 vss 71.2793e-18
c250 n2__i5__net4 vss 71.5683e-18
c251 n42__net4 vss 15.5034e-18
c252 n44__net4 vss 16.4291e-18
c253 n46__net4 vss 12.0074e-18
c254 n38__net4 vss 18.1755e-18
c255 n58__net10 vss 25.2335e-18
c256 n60__net10 vss 22.6563e-18
c257 n62__net10 vss 22.5171e-18
c258 n64__net10 vss 25.7156e-18
c259 n23__rst vss 16.2383e-18
c260 n14__i0__net8 vss 52.1514e-18
c261 n35__rst vss 12.1281e-18
c262 n5__i6__net1 vss 19.0524e-18
c263 n5__i5__net1 vss 17.2551e-18
c264 n4__i0__net11 vss 26.4631e-18
c265 n37__rst vss 11.7846e-18
c266 n7__i7__net1 vss 19.6348e-18
c267 n6__i6__net1 vss 20.6473e-18
c268 n7__i4__net1 vss 20.654e-18
c269 n6__i5__net1 vss 18.6164e-18
c270 n39__rst vss 11.5414e-18
c271 n41__rst vss 11.8142e-18
c272 n7__i0__net10 vss 25.3019e-18
c273 n30__net3 vss 23.5603e-18
c274 n32__net3 vss 22.1025e-18
c275 n34__net3 vss 21.9763e-18
c276 n36__net3 vss 24.7831e-18
c277 n42__rst vss 17.1882e-18
c278 n7__i0__net9 vss 22.004e-18
c279 n3__i7__net2 vss 68.817e-18
c280 n2__i6__net2 vss 72.8273e-18
c281 n3__i4__net2 vss 72.6978e-18
c282 n2__i5__net2 vss 70.283e-18
c283 n13__i0__net8 vss 26.3888e-18
c284 n3__i0__net11 vss 47.3384e-18
c285 n34__net9 vss 25.1404e-18
c286 n36__net9 vss 21.7273e-18
c287 n38__net9 vss 21.5649e-18
c288 n40__net9 vss 24.4437e-18
c289 n14__i0__net1 vss 19.7309e-18
c290 n9__i0__net8 vss 23.2939e-18
c291 n4__i0__i2__net4 vss 22.8263e-18
c292 n6__i0__i3__net4 vss 24.9339e-18
c293 n1__x_out_b_3 vss 23.9143e-18
c294 n4__x_out_b_2 vss 21.8776e-18
c295 n1__x_out_b_1 vss 21.8154e-18
c296 n4__x_out_b_0 vss 20.2559e-18
c297 n5__i0__i3__net5 vss 19.2255e-18
c298 n4__i1__net4 vss 26.9997e-18
c299 n6__i2__net4 vss 23.4371e-18
c300 n4__i3__net4 vss 24.9679e-18
c301 n6__i8__net4 vss 21.8167e-18
c302 n7__i0__i2__net5 vss 20.4407e-18
c303 n6__i0__i3__net5 vss 21.7577e-18
c304 n5__i2__net5 vss 17.3213e-18
c305 n5__i8__net5 vss 15.6984e-18
c306 n7__i1__net5 vss 22.059e-18
c307 n6__i2__net5 vss 21.7179e-18
c308 n7__i3__net5 vss 21.6918e-18
c309 n6__i8__net5 vss 20.0975e-18
c310 n3__i0__i2__net4 vss 75.0121e-18
c311 n2__i0__i3__net4 vss 75.1516e-18
c312 n3__i1__net4 vss 72.9357e-18
c313 n2__i2__net4 vss 75.0074e-18
c314 n3__i3__net4 vss 74.9152e-18
c315 n2__i8__net4 vss 77.2334e-18
c316 n7__clk vss 24.9211e-18
c317 n4__i0__net7 vss 24.4821e-18
c318 n5__i0__i3__net1 vss 20.4802e-18
c319 n10__net10 vss 23.4819e-18
c320 n12__net10 vss 23.3407e-18
c321 n14__net10 vss 23.2074e-18
c322 n16__net10 vss 25.8388e-18
c323 n7__i0__i2__net1 vss 19.4936e-18
c324 n6__i0__i3__net1 vss 19.3631e-18
c325 n5__i2__net1 vss 19.6178e-18
c326 n5__i8__net1 vss 17.9723e-18
c327 n5__rst vss 24.5929e-18
c328 n7__rst vss 23.0364e-18
c329 n7__i1__net1 vss 22.8509e-18
c330 n6__i2__net1 vss 20.7895e-18
c331 n7__i3__net1 vss 20.7939e-18
c332 n6__i8__net1 vss 19.4796e-18
c333 n3__i0__i2__net2 vss 79.0104e-18
c334 n2__i0__i3__net2 vss 77.1314e-18
c335 n2__net3 vss 23.7786e-18
c336 n4__net3 vss 22.1992e-18
c337 n6__net3 vss 22.073e-18
c338 n8__net3 vss 24.3891e-18
c339 n3__i1__net2 vss 76.7795e-18
c340 n2__i2__net2 vss 80.5357e-18
c341 n3__i3__net2 vss 80.4061e-18
c342 n2__i8__net2 vss 85.5464e-18
c343 n2__i0__net3 vss 24.9608e-18
c344 n2__i0__net1 vss 25.8265e-18
c345 n1__clk vss 36.246e-18
c346 n3__rst vss 26.3475e-18
c347 n2__net9 vss 24.7199e-18
c348 n4__net9 vss 25.2594e-18
c349 n6__net9 vss 25.2594e-18
c350 n8__net9 vss 28.0281e-18
c351 n3__y_out_b_3 vss 60.4482e-18
c352 n3__y_out_b_2 vss 61.2402e-18
c353 n3__y_out_b_1 vss 61.2371e-18
c354 n3__y_out_b_0 vss 59.5916e-18
c355 n8__net7 vss 7.80877e-18
c356 n8__net11 vss 7.61985e-18
c357 n5__i7__net4 vss 19.7287e-18
c358 n5__i6__net4 vss 20.7306e-18
c359 n5__i4__net4 vss 20.7269e-18
c360 n5__i5__net4 vss 19.5741e-18
c361 n11__net7 vss 7.80877e-18
c362 n11__net11 vss 7.18244e-18
c363 n4__i7__net5 vss 71.8797e-18
c364 n4__i6__net5 vss 74.8258e-18
c365 n4__i4__net5 vss 75.0262e-18
c366 n4__i5__net5 vss 71.8608e-18
c367 n22__net4 vss 46.4205e-18
c368 n24__net4 vss 46.1507e-18
c369 n26__net4 vss 45.6987e-18
c370 n28__net4 vss 45.4476e-18
c371 n3__net11 vss 117.149e-18
c372 n32__net4 vss 9.55098e-18
c373 n3__net7 vss 8.88971e-18
c374 n35__net4 vss 8.98513e-18
c375 n57__net10 vss 29.9779e-18
c376 n49__net9 vss 25.916e-18
c377 n51__net9 vss 25.916e-18
c378 n59__net10 vss 30.6737e-18
c379 n61__net10 vss 30.669e-18
c380 n53__net9 vss 25.916e-18
c381 n55__net9 vss 25.916e-18
c382 n63__net10 vss 29.9711e-18
c383 n7__i0__net11 vss 30.902e-18
c384 n16__i0__net8 vss 30.6554e-18
c385 n26__rst vss 9.54685e-18
c386 n5__i0__net11 vss 203.95e-18
c387 n4__i7__net1 vss 89.5399e-18
c388 n4__i6__net1 vss 91.9939e-18
c389 n4__i4__net1 vss 91.9845e-18
c390 n4__i5__net1 vss 89.2451e-18
c391 n29__rst vss 6.90627e-18
c392 n6__i0__net10 vss 19.0009e-18
c393 n29__net3 vss 21.5884e-18
c394 n31__net3 vss 22.9014e-18
c395 n33__net3 vss 22.9014e-18
c396 n35__net3 vss 21.2579e-18
c397 n6__i0__net9 vss 19.0685e-18
c398 n3__i0__net9 vss 11.3501e-18
c399 n12__i0__net8 vss 193.877e-18
c400 n11__i0__net8 vss 24.3672e-18
c401 n3__i0__net10 vss 12.6284e-18
c402 n33__net9 vss 30.1314e-18
c403 n41__net10 vss 27.7813e-18
c404 n43__net10 vss 27.7813e-18
c405 n35__net9 vss 30.5009e-18
c406 n37__net9 vss 30.5534e-18
c407 n45__net10 vss 27.7813e-18
c408 n47__net10 vss 27.7813e-18
c409 n39__net9 vss 29.7641e-18
c410 n16__i0__net1 vss 58.226e-18
c411 n8__i0__net8 vss 59.1095e-18
c412 n5__i0__i2__net4 vss 19.5275e-18
c413 n5__i0__i3__net4 vss 20.3194e-18
c414 n3__x_out_b_3 vss 57.9113e-18
c415 n3__x_out_b_2 vss 59.0242e-18
c416 n3__x_out_b_1 vss 59.4831e-18
c417 n3__x_out_b_0 vss 56.6098e-18
c418 n5__i1__net4 vss 19.5209e-18
c419 n5__i2__net4 vss 20.8504e-18
c420 n5__i3__net4 vss 20.8543e-18
c421 n5__i8__net4 vss 19.7892e-18
c422 n4__i0__i2__net5 vss 73.6294e-18
c423 n4__i0__i3__net5 vss 77.1775e-18
c424 n2__i0__net6 vss 43.4881e-18
c425 n4__i0__net6 vss 46.3785e-18
c426 n4__i1__net5 vss 75.6138e-18
c427 n4__i2__net5 vss 77.6539e-18
c428 n4__i3__net5 vss 77.6522e-18
c429 n4__i8__net5 vss 74.894e-18
c430 n2__net4 vss 45.3402e-18
c431 n4__net4 vss 45.044e-18
c432 n6__net4 vss 44.6207e-18
c433 n8__net4 vss 43.8399e-18
c434 n6__clk vss 30.5152e-18
c435 n3__i0__net3 vss 26.8525e-18
c436 n3__i0__net1 vss 26.6537e-18
c437 n3__i0__net7 vss 31.2188e-18
c438 n9__net10 vss 30.0306e-18
c439 n9__net9 vss 26.0082e-18
c440 n11__net9 vss 26.0122e-18
c441 n11__net10 vss 30.6781e-18
c442 n13__net10 vss 30.673e-18
c443 n13__net9 vss 26.0122e-18
c444 n15__net9 vss 26.0122e-18
c445 n15__net10 vss 29.9905e-18
c446 n4__i0__i2__net1 vss 82.4511e-18
c447 n4__i0__i3__net1 vss 87.6707e-18
c448 n4__rst vss 22.0287e-18
c449 n6__rst vss 68.7956e-18
c450 n4__i1__net1 vss 85.6599e-18
c451 n4__i2__net1 vss 88.3338e-18
c452 n4__i3__net1 vss 88.3244e-18
c453 n4__i8__net1 vss 85.3848e-18
c454 n3__net3 vss 22.8113e-18
c455 n5__net3 vss 22.8113e-18
c456 n7__net3 vss 21.1677e-18
c457 n4__clk vss 114.022e-18
c458 n3__net10 vss 29.4931e-18
c459 n3__net9 vss 32.1228e-18
c460 n5__net9 vss 32.1677e-18
c461 n5__net10 vss 29.5632e-18
c462 n7__net10 vss 29.4931e-18
c463 n7__net9 vss 31.3929e-18
c464 n2__clk vss 32.8551e-18
c465 n2__rst vss 33.5597e-18
c466 n220__vdd vss 93.2019e-18
c467 n222__vdd vss 96.3268e-18
c468 n217__vdd vss 7.88231e-18
c469 n218__vdd vss 10.3342e-18
c470 n219__vdd vss 10.3342e-18
c471 n214__vdd vss 11.1587e-18
c472 n215__vdd vss 19.1477e-18
c473 n216__vdd vss 19.1477e-18
c474 n109__net10 vss 669.19e-18
c475 n110__net10 vss 683.664e-18
c476 n111__net10 vss 683.563e-18
c477 n112__net10 vss 608.658e-18
c478 n5__y_out_3 vss 72.8448e-18
c479 n5__y_out_2 vss 71.063e-18
c480 n5__y_out_1 vss 28.0583e-18
c481 n5__y_out_0 vss 28.0675e-18
c482 n39__net7 vss 20.7273e-18
c483 n38__net11 vss 11.9979e-18
c484 n10__y_out_b_3 vss 92.9981e-18
c485 n10__y_out_b_2 vss 92.841e-18
c486 n10__y_out_b_1 vss 63.0101e-18
c487 n10__y_out_b_0 vss 63.0101e-18
c488 n38__net7 vss 46.0824e-18
c489 n37__net11 vss 40.9869e-18
c490 n11__x_out_b_3 vss 722.157e-18
c491 n12__x_out_b_3 vss 103.437e-18
c492 n11__x_out_b_2 vss 102.904e-18
c493 n12__x_out_b_2 vss 722.24e-18
c494 n11__x_out_b_1 vss 722.1e-18
c495 n12__x_out_b_1 vss 103.437e-18
c496 n11__x_out_b_0 vss 102.904e-18
c497 n12__x_out_b_0 vss 722.604e-18
c498 n6__x_out_3 vss 129.244e-18
c499 n7__x_out_3 vss 465.933e-18
c500 n6__x_out_2 vss 465.766e-18
c501 n7__x_out_2 vss 132.416e-18
c502 n6__x_out_1 vss 130.206e-18
c503 n7__x_out_1 vss 465.929e-18
c504 n6__x_out_0 vss 465.766e-18
c505 n7__x_out_0 vss 132.84e-18
c506 n93__net9 vss 584.634e-18
c507 n94__net9 vss 530.717e-18
c508 n95__net9 vss 529.636e-18
c509 n96__net9 vss 484.187e-18
c510 n68__net3 vss 358.568e-18
c511 n69__net3 vss 370.079e-18
c512 n70__net3 vss 369.184e-18
c513 n71__net3 vss 327.106e-18
c514 n37__net7 vss 35.7933e-18
c515 n36__net11 vss 142.368e-18
c516 n64__net3 vss 1.02475e-15
c517 n65__net3 vss 1.02424e-15
c518 n66__net3 vss 1.03891e-15
c519 n67__net3 vss 1.04304e-15
c520 n46__rst vss 358.548e-18
c521 n105__net10 vss 1.10276e-15
c522 n106__net10 vss 1.10235e-15
c523 n107__net10 vss 1.12341e-15
c524 n108__net10 vss 1.123e-15
c525 n89__net9 vss 1.07511e-15
c526 n90__net9 vss 1.07438e-15
c527 n91__net9 vss 1.09713e-15
c528 n92__net9 vss 1.09724e-15
c529 n16__i0__net7 vss 132.334e-18
c530 n1__y_in_3 vss 286.054e-18
c531 n2__y_in_2 vss 295.709e-18
c532 n1__y_in_1 vss 295.59e-18
c533 n2__y_in_0 vss 280.269e-18
c534 n23__i0__net1 vss 102.331e-18
c535 n5__x_out_3 vss 423.867e-18
c536 n5__x_out_2 vss 423.884e-18
c537 n5__x_out_1 vss 423.867e-18
c538 n5__x_out_0 vss 423.884e-18
c539 n10__x_out_b_3 vss 713.811e-18
c540 n9__x_out_b_2 vss 714.015e-18
c541 n10__x_out_b_1 vss 675.174e-18
c542 n9__x_out_b_0 vss 675.221e-18
c543 n21__i0__net1 vss 86.228e-18
c544 n22__i0__net1 vss 246.055e-18
c545 n13__i0__net7 vss 87.7349e-18
c546 n14__i0__net7 vss 241.234e-18
c547 n10__net4 vss 698.682e-18
c548 n11__net4 vss 690.367e-18
c549 n14__net4 vss 677.134e-18
c550 n15__net4 vss 683.438e-18
c551 n7__vdd vss 31.7036e-18
c552 n8__vdd vss 36.0112e-18
c553 n9__vdd vss 36.0112e-18
c554 n25__net3 vss 658.662e-18
c555 n26__net3 vss 660.477e-18
c556 n27__net3 vss 679.757e-18
c557 n28__net3 vss 677.176e-18
c558 n37__net10 vss 241.559e-18
c559 n38__net10 vss 241.223e-18
c560 n39__net10 vss 258.825e-18
c561 n40__net10 vss 258.393e-18
c562 n8__i0__net7 vss 213.301e-18
c563 n29__net9 vss 536.083e-18
c564 n30__net9 vss 535.945e-18
c565 n31__net9 vss 515.475e-18
c566 n32__net9 vss 515.407e-18
c567 n12__i0__net1 vss 280.819e-18
c568 n13__rst vss 476.691e-18
c569 n5__x_in_3 vss 24.5966e-18
c570 n4__x_in_2 vss 25.3626e-18
c571 n5__x_in_1 vss 7.54691e-18
c572 n4__x_in_0 vss 7.37512e-18
c573 n102__net10 vss 47.378e-18
c574 n4__y_out_3 vss 22.6519e-18
c575 n4__y_out_2 vss 21.4416e-18
c576 n4__y_out_1 vss 64.3315e-18
c577 n4__y_out_0 vss 39.7628e-18
c578 n35__net11 vss 40.4686e-18
c579 n9__y_out_b_1 vss 81.4057e-18
c580 n9__y_out_b_0 vss 74.9175e-18
c581 n34__net11 vss 45.8027e-18
c582 n86__net9 vss 116.479e-18
c583 n62__net3 vss 81.7442e-18
c584 n34__net7 vss 16.6489e-18
c585 n32__net11 vss 264.51e-18
c586 n64__net4 vss 132.899e-18
c587 n67__net4 vss 185.405e-18
c588 n68__net4 vss 1.00153e-15
c589 n69__net4 vss 943.712e-18
c590 n70__net4 vss 943.61e-18
c591 n71__net4 vss 963.071e-18
c592 n58__net3 vss 20.0035e-18
c593 n59__net3 vss 511.736e-18
c594 n60__net3 vss 497.092e-18
c595 n61__net3 vss 495.524e-18
c596 n45__rst vss 102.324e-18
c597 n19__i0__net9 vss 136.922e-18
c598 n21__i0__net9 vss 121.358e-18
c599 n19__i0__net10 vss 139.111e-18
c600 n22__i0__net10 vss 206.751e-18
c601 n15__i0__net7 vss 101.719e-18
c602 n8__i0__net11 vss 100.327e-18
c603 n9__i0__net11 vss 108.296e-18
c604 n2__y_in_3 vss 151.435e-18
c605 n1__y_in_2 vss 151.42e-18
c606 n2__y_in_1 vss 49.4358e-18
c607 n1__y_in_0 vss 49.3657e-18
c608 n24__i0__net1 vss 322.548e-18
c609 n25__i0__net1 vss 38.9084e-18
c610 n18__i0__net8 vss 75.1438e-18
c611 n17__i0__net8 vss 359.232e-18
c612 n4__x_out_3 vss 52.7721e-18
c613 n4__x_out_2 vss 54.5441e-18
c614 n4__x_out_1 vss 87.6076e-18
c615 n4__x_out_0 vss 84.822e-18
c616 n9__x_out_b_3 vss 39.5796e-18
c617 n10__x_out_b_2 vss 38.8979e-18
c618 n9__x_out_b_1 vss 78.1851e-18
c619 n10__x_out_b_0 vss 77.4287e-18
c620 n9__net4 vss 641.035e-18
c621 n12__net4 vss 484.908e-18
c622 n13__net4 vss 498.591e-18
c623 n16__net4 vss 525.033e-18
c624 n2__vdd vss 23.3782e-18
c625 n3__vdd vss 23.962e-18
c626 n6__vdd vss 23.962e-18
c627 n21__net3 vss 19.688e-18
c628 n22__net3 vss 19.4164e-18
c629 n23__net3 vss 509.497e-18
c630 n24__net3 vss 508.789e-18
c631 n31__net10 vss 251.593e-18
c632 n35__net10 vss 234.533e-18
c633 n9__i0__net7 vss 114.64e-18
c634 n23__net9 vss 264.313e-18
c635 n27__net9 vss 283.468e-18
c636 n13__i0__net1 vss 108.332e-18
c637 n8__i0__net1 vss 487.385e-18
c638 n9__i0__net1 vss 106.97e-18
c639 n5__i0__net8 vss 155.351e-18
c640 n4__i0__net8 vss 529.052e-18
c641 n8__i0__net6 vss 764.494e-18
c642 n9__i0__net6 vss 780.195e-18
c643 n14__rst vss 442.408e-18
c644 n15__rst vss 277.684e-18
c645 n12__rst vss 25.6961e-18
c646 n4__x_in_1 vss 113.484e-18
c647 n5__x_in_0 vss 113.656e-18
c648 n2__y_out_3 vss 58.3189e-18
c649 n2__y_out_2 vss 58.5855e-18
c650 n2__y_out_1 vss 58.5766e-18
c651 n2__y_out_0 vss 55.899e-18
c652 n80__net9 vss 103.243e-18
c653 n96__net10 vss 29.0799e-18
c654 n32__net7 vss 112.811e-18
c655 n31__net11 vss 70.7506e-18
c656 n6__y_out_b_3 vss 83.8322e-18
c657 n7__y_out_b_2 vss 83.3052e-18
c658 n6__y_out_b_1 vss 32.1943e-18
c659 n7__y_out_b_0 vss 32.223e-18
c660 n77__net9 vss 123.185e-18
c661 n93__net10 vss 46.3411e-18
c662 n13__i7__net4 vss 87.1006e-18
c663 n13__i6__net4 vss 84.8561e-18
c664 n13__i4__net4 vss 84.4378e-18
c665 n13__i5__net4 vss 83.9437e-18
c666 n31__net7 vss 112.867e-18
c667 n30__net11 vss 70.8707e-18
c668 n74__net9 vss 116.816e-18
c669 n90__net10 vss 31.4873e-18
c670 n9__i7__net4 vss 70.6194e-18
c671 n9__i6__net4 vss 69.1321e-18
c672 n9__i4__net4 vss 68.7389e-18
c673 n9__i5__net4 vss 68.6624e-18
c674 n12__i7__net4 vss 107.974e-18
c675 n12__i6__net4 vss 108.545e-18
c676 n12__i4__net4 vss 108.148e-18
c677 n12__i5__net4 vss 108.333e-18
c678 n4__clk_div4_out vss 103.149e-18
c679 n14__i7__net5 vss 140.712e-18
c680 n14__i6__net5 vss 140.514e-18
c681 n14__i4__net5 vss 140.256e-18
c682 n14__i5__net5 vss 139.679e-18
c683 n56__net3 vss 22.4067e-18
c684 n60__net4 vss 109.138e-18
c685 n61__net4 vss 106.125e-18
c686 n62__net4 vss 106.36e-18
c687 n63__net4 vss 108.471e-18
c688 n29__net11 vss 125.625e-18
c689 n59__net4 vss 115.7e-18
c690 n4__clk_div4_out_b vss 136.979e-18
c691 n53__net3 vss 35.2257e-18
c692 n7__i7__net4 vss 146.217e-18
c693 n7__i6__net4 vss 146.149e-18
c694 n7__i4__net4 vss 146.188e-18
c695 n7__i5__net4 vss 145.77e-18
c696 n29__net7 vss 78.2804e-18
c697 n58__net4 vss 118.234e-18
c698 n30__net7 vss 157.917e-18
c699 n11__i7__net5 vss 113.918e-18
c700 n11__i6__net5 vss 112.054e-18
c701 n11__i4__net5 vss 113.266e-18
c702 n11__i5__net5 vss 112.08e-18
c703 n50__net3 vss 50.76e-18
c704 n85__net10 vss 196.592e-18
c705 n69__net9 vss 174.163e-18
c706 n70__net9 vss 173.092e-18
c707 n86__net10 vss 197.001e-18
c708 n87__net10 vss 196.944e-18
c709 n71__net9 vss 174.14e-18
c710 n72__net9 vss 173.092e-18
c711 n88__net10 vss 196.798e-18
c712 n56__net4 vss 118.93e-18
c713 n15__i0__net11 vss 137.629e-18
c714 n17__i0__net10 vss 150.732e-18
c715 n25__i0__net8 vss 237.692e-18
c716 n44__rst vss 129.042e-18
c717 n12__i7__net2 vss 200.348e-18
c718 n12__i6__net2 vss 200.272e-18
c719 n12__i4__net2 vss 200.284e-18
c720 n12__i5__net2 vss 200.291e-18
c721 n53__net4 vss 134.932e-18
c722 n14__i0__net11 vss 229.691e-18
c723 n43__rst vss 143.574e-18
c724 n15__i0__net10 vss 88.7786e-18
c725 n16__i7__net1 vss 111.497e-18
c726 n16__i6__net1 vss 111.285e-18
c727 n16__i4__net1 vss 111.036e-18
c728 n16__i5__net1 vss 111.172e-18
c729 n50__net4 vss 110.427e-18
c730 n38__net3 vss 496.332e-18
c731 n17__i0__net9 vss 251.613e-18
c732 n14__i7__net1 vss 251.394e-18
c733 n14__i6__net1 vss 251.068e-18
c734 n14__i4__net1 vss 251.332e-18
c735 n14__i5__net1 vss 251.068e-18
c736 n10__i0__net10 vss 170.875e-18
c737 n61__net9 vss 320.398e-18
c738 n63__net9 vss 320.495e-18
c739 n65__net9 vss 320.445e-18
c740 n67__net9 vss 320.173e-18
c741 n12__i0__net9 vss 54.2819e-18
c742 n77__net10 vss 279.862e-18
c743 n78__net10 vss 251.063e-18
c744 n79__net10 vss 250.849e-18
c745 n80__net10 vss 281.78e-18
c746 n81__net10 vss 281.588e-18
c747 n82__net10 vss 230.347e-18
c748 n83__net10 vss 230.194e-18
c749 n84__net10 vss 280.754e-18
c750 n28__net7 vss 270.608e-18
c751 n24__i0__net8 vss 293.404e-18
c752 n11__i0__net9 vss 71.5518e-18
c753 n62__net9 vss 283.944e-18
c754 n64__net9 vss 283.84e-18
c755 n66__net9 vss 260.973e-18
c756 n68__net9 vss 260.344e-18
c757 n13__i0__net11 vss 99.0114e-18
c758 n28__net11 vss 209.874e-18
c759 n9__i0__net9 vss 138.03e-18
c760 n4__i7__net2 vss 231.967e-18
c761 n4__i6__net2 vss 232.156e-18
c762 n4__i4__net2 vss 232.156e-18
c763 n4__i5__net2 vss 231.777e-18
c764 n23__i0__net8 vss 118.46e-18
c765 n8__i0__net10 vss 71.6768e-18
c766 n11__i7__net1 vss 240.696e-18
c767 n11__i6__net1 vss 240.26e-18
c768 n11__i4__net1 vss 240.408e-18
c769 n11__i5__net1 vss 240.26e-18
c770 n66__net10 vss 146.448e-18
c771 n70__net10 vss 178.661e-18
c772 n72__net10 vss 146.393e-18
c773 n76__net10 vss 178.661e-18
c774 n18__i0__net7 vss 47.3095e-18
c775 n11__i0__net11 vss 44.8734e-18
c776 n57__net9 vss 252.98e-18
c777 n58__net9 vss 250.993e-18
c778 n59__net9 vss 251.898e-18
c779 n60__net9 vss 251.069e-18
c780 n4__y_in_3 vss 89.5842e-18
c781 n4__y_in_2 vss 88.4117e-18
c782 n4__y_in_1 vss 190.451e-18
c783 n4__y_in_0 vss 190.466e-18
c784 n27__i0__net1 vss 51.5957e-18
c785 n21__i0__net8 vss 32.1284e-18
c786 n2__x_out_3 vss 80.2436e-18
c787 n2__x_out_2 vss 79.5742e-18
c788 n2__x_out_1 vss 45.1064e-18
c789 n2__x_out_0 vss 45.0614e-18
c790 n13__i0__i2__net4 vss 94.9799e-18
c791 n13__i0__i3__net4 vss 94.9728e-18
c792 n6__x_out_b_3 vss 43.7112e-18
c793 n7__x_out_b_2 vss 43.5285e-18
c794 n6__x_out_b_1 vss 43.5285e-18
c795 n7__x_out_b_0 vss 43.5693e-18
c796 n9__i0__i2__net4 vss 73.5744e-18
c797 n9__i0__i3__net4 vss 77.5414e-18
c798 n12__i0__i2__net4 vss 111.674e-18
c799 n12__i0__i3__net4 vss 112.452e-18
c800 n13__i1__net4 vss 87.742e-18
c801 n13__i2__net4 vss 88.493e-18
c802 n13__i3__net4 vss 85.3142e-18
c803 n13__i8__net4 vss 86.1544e-18
c804 n14__i0__i2__net5 vss 140.036e-18
c805 n14__i0__i3__net5 vss 140.453e-18
c806 n9__i1__net4 vss 73.0645e-18
c807 n9__i2__net4 vss 75.2035e-18
c808 n9__i3__net4 vss 72.9342e-18
c809 n9__i8__net4 vss 72.5514e-18
c810 n12__i1__net4 vss 112.289e-18
c811 n12__i2__net4 vss 112.201e-18
c812 n12__i3__net4 vss 112.364e-18
c813 n12__i8__net4 vss 112.132e-18
c814 n10__i0__net6 vss 456.556e-18
c815 n11__i0__net6 vss 452.524e-18
c816 n14__i1__net5 vss 135.83e-18
c817 n14__i2__net5 vss 136.11e-18
c818 n14__i3__net5 vss 135.389e-18
c819 n14__i8__net5 vss 136.156e-18
c820 n17__net4 vss 70.9517e-18
c821 n18__net4 vss 70.9358e-18
c822 n19__net4 vss 71.3495e-18
c823 n20__net4 vss 68.594e-18
c824 n7__i0__i2__net4 vss 148.747e-18
c825 n7__i0__i3__net4 vss 150.889e-18
c826 n11__i0__i2__net5 vss 116.384e-18
c827 n11__i0__i3__net5 vss 113.735e-18
c828 n1__vdd vss 142.932e-18
c829 n4__vdd vss 235.605e-18
c830 n5__vdd vss 236.173e-18
c831 n7__i1__net4 vss 170.261e-18
c832 n7__i2__net4 vss 170.354e-18
c833 n7__i3__net4 vss 170.352e-18
c834 n7__i8__net4 vss 170.182e-18
c835 n18__clk vss 198.364e-18
c836 n11__i0__net3 vss 186.572e-18
c837 n20__i0__net1 vss 186.504e-18
c838 n12__i0__net7 vss 195.402e-18
c839 n11__i1__net5 vss 117.209e-18
c840 n11__i2__net5 vss 117.779e-18
c841 n11__i3__net5 vss 117.398e-18
c842 n11__i8__net5 vss 117.894e-18
c843 n53__net10 vss 192.35e-18
c844 n45__net9 vss 167.303e-18
c845 n46__net9 vss 167.199e-18
c846 n54__net10 vss 192.286e-18
c847 n55__net10 vss 192.124e-18
c848 n47__net9 vss 167.239e-18
c849 n48__net9 vss 167.199e-18
c850 n56__net10 vss 192.335e-18
c851 n5__i0__i2__net2 vss 204.405e-18
c852 n5__i0__i3__net2 vss 206.499e-18
c853 n16__i0__i2__net1 vss 106.538e-18
c854 n16__i0__i3__net1 vss 111.874e-18
c855 n5__i1__net2 vss 206.673e-18
c856 n5__i2__net2 vss 206.676e-18
c857 n5__i3__net2 vss 206.673e-18
c858 n5__i8__net2 vss 206.671e-18
c859 n17__rst vss 371.7e-18
c860 n19__rst vss 221.033e-18
c861 n14__i0__i2__net1 vss 252.537e-18
c862 n14__i0__i3__net1 vss 251.261e-18
c863 n10__i0__net3 vss 322.42e-18
c864 n19__i0__net1 vss 322.724e-18
c865 n16__i1__net1 vss 111.864e-18
c866 n16__i2__net1 vss 112.071e-18
c867 n16__i3__net1 vss 111.673e-18
c868 n16__i8__net1 vss 111.958e-18
c869 n15__clk vss 273.307e-18
c870 n16__clk vss 217.53e-18
c871 n10__i0__net7 vss 183.252e-18
c872 n11__i0__net7 vss 284.325e-18
c873 n10__net3 vss 509.593e-18
c874 n12__net3 vss 508.66e-18
c875 n14__i1__net1 vss 253.644e-18
c876 n14__i2__net1 vss 253.121e-18
c877 n14__i3__net1 vss 253.508e-18
c878 n14__i8__net1 vss 253.128e-18
c879 n9__i0__net3 vss 266.729e-18
c880 n18__i0__net1 vss 254.156e-18
c881 n41__net9 vss 320.702e-18
c882 n42__net9 vss 320.082e-18
c883 n43__net9 vss 320.488e-18
c884 n44__net9 vss 319.911e-18
c885 n49__net10 vss 281.954e-18
c886 n29__net10 vss 251.275e-18
c887 n50__net10 vss 281.872e-18
c888 n51__net10 vss 282.28e-18
c889 n33__net10 vss 233.774e-18
c890 n52__net10 vss 281.017e-18
c891 n4__i0__i2__net2 vss 236.069e-18
c892 n4__i0__i3__net2 vss 238.071e-18
c893 n21__net9 vss 264.443e-18
c894 n25__net9 vss 284.782e-18
c895 n11__i0__i2__net1 vss 235.001e-18
c896 n11__i0__i3__net1 vss 240.636e-18
c897 n13__clk vss 65.9282e-18
c898 n7__i0__net7 vss 88.2895e-18
c899 n4__i1__net2 vss 238.737e-18
c900 n4__i2__net2 vss 238.802e-18
c901 n4__i3__net2 vss 238.756e-18
c902 n4__i8__net2 vss 238.7e-18
c903 n8__i0__net3 vss 235.266e-18
c904 n10__i0__net1 vss 159.469e-18
c905 n6__i0__net1 vss 138.883e-18
c906 n2__i0__net8 vss 126.337e-18
c907 n11__i1__net1 vss 237.027e-18
c908 n11__i2__net1 vss 236.543e-18
c909 n11__i3__net1 vss 236.86e-18
c910 n11__i8__net1 vss 236.693e-18
c911 n6__i0__net3 vss 135.652e-18
c912 n6__i0__net6 vss 109.944e-18
c913 n18__net10 vss 177.921e-18
c914 n22__net10 vss 176.865e-18
c915 n24__net10 vss 177.841e-18
c916 n28__net10 vss 176.971e-18
c917 n17__net9 vss 253.554e-18
c918 n18__net9 vss 252.209e-18
c919 n19__net9 vss 253.08e-18
c920 n20__net9 vss 252.428e-18
c921 n8__clk vss 51.3678e-18
c922 n2__x_in_3 vss 174.678e-18
c923 n2__x_in_2 vss 173.497e-18
c924 n2__x_in_1 vss 77.9716e-18
c925 n2__x_in_0 vss 77.9491e-18
c926 n16__vdd vss 6.36068e-15
c927 n97__vdd vss 1.55157e-15
c928 n157__vdd vss 1.55127e-15
c929 n13__vdd vss 60.8322e-18
c930 n26__vdd vss 52.9428e-18
c931 n3__y_out_3 vss 79.0014e-18
c932 n1__y_out_2 vss 78.7792e-18
c933 n3__y_out_1 vss 79.0014e-18
c934 n1__y_out_0 vss 80.6081e-18
c935 n81__net9 vss 66.2902e-18
c936 n95__net10 vss 112.118e-18
c937 n94__vdd vss 87.587e-18
c938 n114__vdd vss 87.8192e-18
c939 n154__vdd vss 87.587e-18
c940 n174__vdd vss 88.1537e-18
c941 n28__vdd vss 106.33e-18
c942 n27__vdd vss 99.7941e-18
c943 n7__y_out_b_3 vss 55.5805e-18
c944 n8__y_out_b_2 vss 55.6321e-18
c945 n7__y_out_b_1 vss 55.6321e-18
c946 n8__y_out_b_0 vss 55.642e-18
c947 n78__net9 vss 66.1035e-18
c948 n92__net10 vss 117.526e-18
c949 n116__vdd vss 63.1585e-18
c950 n115__vdd vss 63.0297e-18
c951 n176__vdd vss 63.009e-18
c952 n175__vdd vss 63.1081e-18
c953 n30__vdd vss 106.319e-18
c954 n29__vdd vss 100.258e-18
c955 n118__vdd vss 56.8539e-18
c956 n117__vdd vss 56.8792e-18
c957 n178__vdd vss 56.8792e-18
c958 n177__vdd vss 56.9201e-18
c959 n75__net9 vss 65.631e-18
c960 n89__net10 vss 113.969e-18
c961 n10__i7__net4 vss 44.785e-18
c962 n10__i6__net4 vss 44.6717e-18
c963 n10__i4__net4 vss 44.7641e-18
c964 n10__i5__net4 vss 44.6813e-18
c965 n32__vdd vss 87.6598e-18
c966 n31__vdd vss 49.1619e-18
c967 n120__vdd vss 89.6768e-18
c968 n119__vdd vss 89.786e-18
c969 n180__vdd vss 89.6713e-18
c970 n179__vdd vss 89.7974e-18
c971 n33__vdd vss 50.5464e-18
c972 n2__clk_div4_out vss 51.7072e-18
c973 n15__i7__net5 vss 831.967e-21
c974 n15__i6__net5 vss 827.251e-21
c975 n15__i4__net5 vss 847.984e-21
c976 n15__i5__net5 vss 900.802e-21
c977 n55__net3 vss 113.503e-18
c978 n34__vdd vss 105.475e-18
c979 n122__vdd vss 26.573e-18
c980 n121__vdd vss 26.3812e-18
c981 n182__vdd vss 26.3897e-18
c982 n181__vdd vss 25.7351e-18
c983 n35__vdd vss 99.8201e-18
c984 n1__clk_div4_out_b vss 150.359e-18
c985 n52__net3 vss 123.326e-18
c986 n124__vdd vss 50.7945e-18
c987 n123__vdd vss 51.2323e-18
c988 n184__vdd vss 51.1505e-18
c989 n183__vdd vss 50.6981e-18
c990 n36__vdd vss 61.8098e-18
c991 n37__vdd vss 96.4096e-18
c992 n9__i7__net5 vss 39.4895e-18
c993 n9__i6__net5 vss 37.261e-18
c994 n9__i4__net5 vss 39.496e-18
c995 n9__i5__net5 vss 37.261e-18
c996 n49__net3 vss 121.863e-18
c997 n12__i7__net5 vss 83.2328e-18
c998 n13__i6__net5 vss 83.2569e-18
c999 n12__i4__net5 vss 83.0991e-18
c1000 n13__i5__net5 vss 83.2569e-18
c1001 n38__vdd vss 78.3423e-18
c1002 n44__vdd vss 62.8597e-18
c1003 n10__i7__net2 vss 80.5716e-18
c1004 n5__i6__net2 vss 80.3863e-18
c1005 n10__i4__net2 vss 80.5716e-18
c1006 n5__i5__net2 vss 80.3863e-18
c1007 n57__net4 vss 67.6393e-18
c1008 n126__vdd vss 90.4205e-18
c1009 n125__vdd vss 90.4714e-18
c1010 n186__vdd vss 90.4193e-18
c1011 n185__vdd vss 90.4702e-18
c1012 n16__i0__net10 vss 66.0976e-18
c1013 n45__vdd vss 105.497e-18
c1014 n8__i7__net2 vss 47.234e-18
c1015 n10__i6__net2 vss 47.121e-18
c1016 n8__i4__net2 vss 47.2348e-18
c1017 n10__i5__net2 vss 47.1218e-18
c1018 n41__vdd vss 135.502e-18
c1019 n54__net4 vss 66.947e-18
c1020 n128__vdd vss 94.6127e-18
c1021 n127__vdd vss 94.59e-18
c1022 n188__vdd vss 94.6144e-18
c1023 n187__vdd vss 94.5917e-18
c1024 n51__vdd vss 107.34e-18
c1025 n47__vdd vss 136.723e-18
c1026 n51__net4 vss 66.3758e-18
c1027 n16__i0__net9 vss 108.814e-18
c1028 n52__vdd vss 81.1368e-18
c1029 n9__i0__net10 vss 84.8376e-18
c1030 n50__vdd vss 112.036e-18
c1031 n25__net7 vss 116.32e-18
c1032 n58__vdd vss 77.0179e-18
c1033 n55__vdd vss 114.628e-18
c1034 n130__vdd vss 90.6236e-18
c1035 n129__vdd vss 90.6738e-18
c1036 n190__vdd vss 90.6738e-18
c1037 n189__vdd vss 90.0242e-18
c1038 n8__i0__net9 vss 79.1945e-18
c1039 n26__net11 vss 48.7254e-18
c1040 n63__vdd vss 88.4017e-18
c1041 n9__i7__net1 vss 39.6551e-18
c1042 n9__i6__net1 vss 37.2963e-18
c1043 n9__i4__net1 vss 39.6551e-18
c1044 n9__i5__net1 vss 37.2963e-18
c1045 n12__i7__net1 vss 86.5651e-18
c1046 n13__i6__net1 vss 86.5975e-18
c1047 n12__i4__net1 vss 86.5651e-18
c1048 n13__i5__net1 vss 86.5975e-18
c1049 n19__i0__net7 vss 84.1005e-18
c1050 n10__i0__net11 vss 91.8674e-18
c1051 n5__y_in_3 vss 49.6299e-18
c1052 n3__y_in_2 vss 49.4623e-18
c1053 n5__y_in_1 vss 49.6621e-18
c1054 n3__y_in_0 vss 49.4623e-18
c1055 n66__vdd vss 85.3509e-18
c1056 n62__vdd vss 87.7637e-18
c1057 n28__i0__net1 vss 53.3861e-18
c1058 n22__i0__net8 vss 55.574e-18
c1059 n3__x_out_3 vss 94.0231e-18
c1060 n1__x_out_2 vss 93.7775e-18
c1061 n3__x_out_1 vss 94.0231e-18
c1062 n1__x_out_0 vss 93.7775e-18
c1063 n69__vdd vss 64.3271e-18
c1064 n65__vdd vss 68.358e-18
c1065 n132__vdd vss 91.8746e-18
c1066 n131__vdd vss 91.8746e-18
c1067 n192__vdd vss 91.8746e-18
c1068 n191__vdd vss 91.8746e-18
c1069 n72__vdd vss 57.6707e-18
c1070 n68__vdd vss 59.3292e-18
c1071 n7__x_out_b_3 vss 55.9984e-18
c1072 n8__x_out_b_2 vss 56.0177e-18
c1073 n7__x_out_b_1 vss 56.0177e-18
c1074 n8__x_out_b_0 vss 56.0177e-18
c1075 n10__i0__i2__net4 vss 44.0446e-18
c1076 n10__i0__i3__net4 vss 42.9606e-18
c1077 n134__vdd vss 63.0628e-18
c1078 n133__vdd vss 62.9982e-18
c1079 n194__vdd vss 62.9982e-18
c1080 n193__vdd vss 62.9982e-18
c1081 n75__vdd vss 89.5323e-18
c1082 n71__vdd vss 91.7198e-18
c1083 n136__vdd vss 56.9525e-18
c1084 n135__vdd vss 56.9779e-18
c1085 n196__vdd vss 56.9779e-18
c1086 n195__vdd vss 56.9525e-18
c1087 n10__i1__net4 vss 45.1433e-18
c1088 n10__i2__net4 vss 44.989e-18
c1089 n10__i3__net4 vss 45.107e-18
c1090 n10__i8__net4 vss 44.989e-18
c1091 n78__vdd vss 26.2735e-18
c1092 n74__vdd vss 26.2967e-18
c1093 n138__vdd vss 89.7842e-18
c1094 n137__vdd vss 89.5671e-18
c1095 n198__vdd vss 89.7965e-18
c1096 n197__vdd vss 89.5671e-18
c1097 n82__vdd vss 50.0529e-18
c1098 n77__vdd vss 49.4138e-18
c1099 n140__vdd vss 25.4994e-18
c1100 n139__vdd vss 25.1057e-18
c1101 n200__vdd vss 25.3773e-18
c1102 n199__vdd vss 24.666e-18
c1103 n9__i0__i2__net5 vss 39.3832e-18
c1104 n9__i0__i3__net5 vss 37.0994e-18
c1105 n144__vdd vss 48.791e-18
c1106 n141__vdd vss 49.4901e-18
c1107 n204__vdd vss 49.4901e-18
c1108 n201__vdd vss 49.0115e-18
c1109 n12__i0__i2__net5 vss 82.5608e-18
c1110 n13__i0__i3__net5 vss 84.6139e-18
c1111 n11__i0__i2__net2 vss 79.2827e-18
c1112 n6__i0__i3__net2 vss 79.2827e-18
c1113 n9__i1__net5 vss 40.9353e-18
c1114 n9__i2__net5 vss 38.5583e-18
c1115 n9__i3__net5 vss 40.9328e-18
c1116 n9__i8__net5 vss 38.5583e-18
c1117 n85__vdd vss 90.2119e-18
c1118 n81__vdd vss 91.0166e-18
c1119 n12__i1__net5 vss 82.7199e-18
c1120 n13__i2__net5 vss 82.8057e-18
c1121 n12__i3__net5 vss 82.7732e-18
c1122 n13__i8__net5 vss 82.8057e-18
c1123 n9__i0__i2__net2 vss 46.5818e-18
c1124 n11__i0__i3__net2 vss 46.5027e-18
c1125 n11__i1__net2 vss 79.6987e-18
c1126 n6__i2__net2 vss 79.4835e-18
c1127 n11__i3__net2 vss 79.6987e-18
c1128 n6__i8__net2 vss 79.4835e-18
c1129 n88__vdd vss 94.8013e-18
c1130 n84__vdd vss 94.9601e-18
c1131 n147__vdd vss 89.5375e-18
c1132 n143__vdd vss 89.7468e-18
c1133 n207__vdd vss 89.5467e-18
c1134 n203__vdd vss 89.7468e-18
c1135 n9__i1__net2 vss 47.0102e-18
c1136 n11__i2__net2 vss 46.8972e-18
c1137 n9__i3__net2 vss 47.0102e-18
c1138 n11__i8__net2 vss 46.8972e-18
c1139 n151__vdd vss 94.8893e-18
c1140 n146__vdd vss 94.8893e-18
c1141 n211__vdd vss 94.8893e-18
c1142 n206__vdd vss 94.8893e-18
c1143 n92__vdd vss 91.7886e-18
c1144 n87__vdd vss 90.6807e-18
c1145 n9__i0__i2__net1 vss 39.9621e-18
c1146 n9__i0__i3__net1 vss 37.0328e-18
c1147 n153__vdd vss 91.9347e-18
c1148 n150__vdd vss 92.1307e-18
c1149 n213__vdd vss 92.1307e-18
c1150 n210__vdd vss 91.6474e-18
c1151 n12__i0__i2__net1 vss 87.13e-18
c1152 n13__i0__i3__net1 vss 86.2857e-18
c1153 n7__i0__net1 vss 57.7295e-18
c1154 n9__i1__net1 vss 40.5958e-18
c1155 n9__i2__net1 vss 38.3284e-18
c1156 n9__i3__net1 vss 40.6761e-18
c1157 n9__i8__net1 vss 38.3161e-18
c1158 n7__i0__net3 vss 78.7391e-18
c1159 n5__i0__net6 vss 91.0422e-18
c1160 n12__i1__net1 vss 86.7815e-18
c1161 n13__i2__net1 vss 86.819e-18
c1162 n12__i3__net1 vss 86.7868e-18
c1163 n13__i8__net1 vss 86.819e-18
c1164 n93__vdd vss 45.1172e-18
c1165 n91__vdd vss 36.7852e-18
c1166 n3__x_in_3 vss 53.5993e-18
c1167 n1__x_in_2 vss 53.4084e-18
c1168 n3__x_in_1 vss 53.5993e-18
c1169 n1__x_in_0 vss 53.4084e-18
c1170 n1__y_out_3 vss 42.8067e-18
c1171 n3__y_out_2 vss 48.6596e-18
c1172 n1__y_out_1 vss 48.5637e-18
c1173 n3__y_out_0 vss 46.8861e-18
c1174 n79__net9 vss 75.0354e-18
c1175 n97__net10 vss 77.7968e-18
c1176 n8__y_out_b_3 vss 51.5596e-18
c1177 n6__y_out_b_2 vss 49.0099e-18
c1178 n8__y_out_b_1 vss 49.0099e-18
c1179 n6__y_out_b_0 vss 47.4597e-18
c1180 n76__net9 vss 78.6917e-18
c1181 n94__net10 vss 86.1873e-18
c1182 n73__net9 vss 77.4497e-18
c1183 n91__net10 vss 79.4947e-18
c1184 n8__i7__net4 vss 61.3326e-18
c1185 n8__i6__net4 vss 61.3269e-18
c1186 n8__i4__net4 vss 61.3269e-18
c1187 n8__i5__net4 vss 58.2525e-18
c1188 n1__clk_div4_out vss 89.1751e-18
c1189 n57__net3 vss 77.0714e-18
c1190 n54__net3 vss 88.506e-18
c1191 n8__i7__net5 vss 35.1184e-18
c1192 n8__i6__net5 vss 36.1874e-18
c1193 n8__i4__net5 vss 33.9302e-18
c1194 n8__i5__net5 vss 36.3786e-18
c1195 n51__net3 vss 81.2491e-18
c1196 n13__i7__net5 vss 56.1541e-18
c1197 n12__i6__net5 vss 54.218e-18
c1198 n13__i4__net5 vss 54.2967e-18
c1199 n12__i5__net5 vss 54.5858e-18
c1200 n5__i7__net2 vss 33.7749e-18
c1201 n9__i6__net2 vss 34.1049e-18
c1202 n5__i4__net2 vss 34.0185e-18
c1203 n9__i5__net2 vss 33.0767e-18
c1204 n55__net4 vss 76.3858e-18
c1205 n18__i0__net10 vss 46.6151e-18
c1206 n11__i7__net2 vss 57.1946e-18
c1207 n8__i6__net2 vss 56.979e-18
c1208 n11__i4__net2 vss 57.007e-18
c1209 n8__i5__net2 vss 57.0639e-18
c1210 n43__vdd vss 90.3585e-18
c1211 n52__net4 vss 78.6864e-18
c1212 n49__net4 vss 78.203e-18
c1213 n18__i0__net9 vss 50.5204e-18
c1214 n15__i7__net1 vss 63.7027e-18
c1215 n15__i6__net1 vss 63.4971e-18
c1216 n15__i4__net1 vss 63.478e-18
c1217 n15__i5__net1 vss 62.0367e-18
c1218 n11__i0__net10 vss 72.0213e-18
c1219 n57__vdd vss 102.544e-18
c1220 n10__i0__net9 vss 28.8459e-18
c1221 n25__net11 vss 110.155e-18
c1222 n8__i7__net1 vss 34.9644e-18
c1223 n8__i6__net1 vss 35.1831e-18
c1224 n8__i4__net1 vss 33.0671e-18
c1225 n8__i5__net1 vss 34.4648e-18
c1226 n13__i7__net1 vss 56.7878e-18
c1227 n12__i6__net1 vss 55.2084e-18
c1228 n13__i4__net1 vss 55.2586e-18
c1229 n12__i5__net1 vss 55.3402e-18
c1230 n17__i0__net7 vss 49.3654e-18
c1231 n12__i0__net11 vss 48.5664e-18
c1232 n3__y_in_3 vss 55.9187e-18
c1233 n5__y_in_2 vss 56.0338e-18
c1234 n3__y_in_1 vss 55.9077e-18
c1235 n5__y_in_0 vss 55.6026e-18
c1236 n29__i0__net1 vss 46.7044e-18
c1237 n20__i0__net8 vss 46.8828e-18
c1238 n1__x_out_3 vss 55.5582e-18
c1239 n3__x_out_2 vss 54.3476e-18
c1240 n1__x_out_1 vss 54.2391e-18
c1241 n3__x_out_0 vss 53.3582e-18
c1242 n8__x_out_b_3 vss 55.7929e-18
c1243 n6__x_out_b_2 vss 51.4121e-18
c1244 n8__x_out_b_1 vss 51.4121e-18
c1245 n6__x_out_b_0 vss 52.5341e-18
c1246 n8__i0__i2__net4 vss 61.0557e-18
c1247 n8__i0__i3__net4 vss 62.9968e-18
c1248 n8__i1__net4 vss 62.157e-18
c1249 n8__i2__net4 vss 60.9892e-18
c1250 n8__i3__net4 vss 60.9892e-18
c1251 n8__i8__net4 vss 61.6746e-18
c1252 n8__i0__i2__net5 vss 34.7004e-18
c1253 n8__i0__i3__net5 vss 36.5699e-18
c1254 n13__i0__i2__net5 vss 54.2751e-18
c1255 n12__i0__i3__net5 vss 54.365e-18
c1256 n6__i0__i2__net2 vss 32.6754e-18
c1257 n10__i0__i3__net2 vss 33.6148e-18
c1258 n8__i1__net5 vss 32.4811e-18
c1259 n8__i2__net5 vss 34.6642e-18
c1260 n8__i3__net5 vss 32.4785e-18
c1261 n8__i8__net5 vss 35.4478e-18
c1262 n13__i1__net5 vss 53.3295e-18
c1263 n12__i2__net5 vss 53.1403e-18
c1264 n13__i3__net5 vss 52.6768e-18
c1265 n12__i8__net5 vss 53.9942e-18
c1266 n12__i0__i2__net2 vss 58.7667e-18
c1267 n9__i0__i3__net2 vss 59.7657e-18
c1268 n6__i1__net2 vss 32.643e-18
c1269 n10__i2__net2 vss 32.5289e-18
c1270 n6__i3__net2 vss 32.4336e-18
c1271 n10__i8__net2 vss 33.2217e-18
c1272 n12__i1__net2 vss 59.1328e-18
c1273 n9__i2__net2 vss 58.3282e-18
c1274 n12__i3__net2 vss 58.3527e-18
c1275 n9__i8__net2 vss 58.9094e-18
c1276 n15__i0__i2__net1 vss 62.0426e-18
c1277 n15__i0__i3__net1 vss 62.6659e-18
c1278 n15__i1__net1 vss 63.8327e-18
c1279 n15__i2__net1 vss 63.2224e-18
c1280 n15__i3__net1 vss 63.2032e-18
c1281 n15__i8__net1 vss 63.5334e-18
c1282 n8__i0__i2__net1 vss 33.5086e-18
c1283 n8__i0__i3__net1 vss 36.4805e-18
c1284 n13__i0__i2__net1 vss 55.7372e-18
c1285 n12__i0__i3__net1 vss 56.4951e-18
c1286 n5__i0__net1 vss 57.5718e-18
c1287 n3__i0__net8 vss 63.1345e-18
c1288 n8__i1__net1 vss 33.1876e-18
c1289 n8__i2__net1 vss 34.8656e-18
c1290 n8__i3__net1 vss 32.775e-18
c1291 n8__i8__net1 vss 36.34e-18
c1292 n5__i0__net3 vss 58.1735e-18
c1293 n7__i0__net6 vss 38.2584e-18
c1294 n13__i1__net1 vss 56.8506e-18
c1295 n12__i2__net1 vss 56.8982e-18
c1296 n13__i3__net1 vss 56.912e-18
c1297 n12__i8__net1 vss 57.4999e-18
c1298 n1__x_in_3 vss 49.5957e-18
c1299 n3__x_in_2 vss 49.2134e-18
c1300 n1__x_in_1 vss 49.0561e-18
c1301 n3__x_in_0 vss 50.5215e-18
c1302 n2__i1__net1 vss 16.8064e-18
c1303 n3__i1__net1 vss 8.85348e-18
c1304 n2__i2__net1 vss 16.4865e-18
c1305 n3__i2__net1 vss 8.84604e-18
c1306 n2__i3__net1 vss 16.8035e-18
c1307 n3__i3__net1 vss 9.19344e-18
c1308 n2__i8__net1 vss 15.4046e-18
c1309 n3__i8__net1 vss 7.81321e-18
c1310 n2__i0__i2__net1 vss 16.2745e-18
c1311 n3__i0__i2__net1 vss 8.12086e-18
c1312 n2__i0__i3__net1 vss 15.7722e-18
c1313 n3__i0__i3__net1 vss 8.30894e-18
c1314 n2__i1__net5 vss 16.8615e-18
c1315 n3__i1__net5 vss 10.5627e-18
c1316 n2__i2__net5 vss 19.0843e-18
c1317 n3__i2__net5 vss 10.2793e-18
c1318 n2__i3__net5 vss 17.694e-18
c1319 n3__i3__net5 vss 10.6226e-18
c1320 n2__i8__net5 vss 18.0938e-18
c1321 n3__i8__net5 vss 9.28465e-18
c1322 n9__clk vss 27.2648e-18
c1323 n10__clk vss 34.5409e-18
c1324 n9__rst vss 17.8635e-18
c1325 n10__rst vss 33.5748e-18
c1326 n2__i0__i2__net5 vss 18.0268e-18
c1327 n3__i0__i2__net5 vss 8.93933e-18
c1328 n2__i0__i3__net5 vss 17.588e-18
c1329 n3__i0__i3__net5 vss 9.25057e-18
c1330 n19__net10 vss 53.7153e-18
c1331 n20__net10 vss 53.8725e-18
c1332 n25__net10 vss 53.7217e-18
c1333 n26__net10 vss 53.8725e-18
c1334 n2__x_out_b_3 vss 9.56972e-18
c1335 n2__x_out_b_2 vss 10.1258e-18
c1336 n2__x_out_b_1 vss 9.54338e-18
c1337 n2__x_out_b_0 vss 10.1258e-18
c1338 n6__i0__net7 vss 33.6468e-18
c1339 n15__i0__net1 vss 11.166e-18
c1340 n7__i0__net8 vss 9.11932e-18
c1341 n2__i0__net10 vss 10.7723e-18
c1342 n9__net3 vss 45.6161e-18
c1343 n11__net3 vss 43.1337e-18
c1344 n13__net3 vss 44.2171e-18
c1345 n14__net3 vss 45.3372e-18
c1346 n15__net3 vss 45.6161e-18
c1347 n17__net3 vss 43.9352e-18
c1348 n19__net3 vss 43.2688e-18
c1349 n20__net3 vss 45.3372e-18
c1350 n2__i0__net9 vss 11.3653e-18
c1351 n7__i1__net2 vss 89.4041e-18
c1352 n8__i1__net2 vss 57.7263e-18
c1353 n7__i2__net2 vss 88.8825e-18
c1354 n8__i2__net2 vss 57.2045e-18
c1355 n7__i3__net2 vss 88.3159e-18
c1356 n8__i3__net2 vss 57.5145e-18
c1357 n7__i8__net2 vss 88.8591e-18
c1358 n8__i8__net2 vss 56.775e-18
c1359 n2__i7__net1 vss 17.2096e-18
c1360 n3__i7__net1 vss 9.4067e-18
c1361 n2__i6__net1 vss 16.9032e-18
c1362 n3__i6__net1 vss 8.8989e-18
c1363 n2__i4__net1 vss 17.2204e-18
c1364 n3__i4__net1 vss 9.2441e-18
c1365 n2__i5__net1 vss 15.8187e-18
c1366 n3__i5__net1 vss 7.92248e-18
c1367 n7__i0__i2__net2 vss 88.351e-18
c1368 n8__i0__i2__net2 vss 54.4369e-18
c1369 n7__i0__i3__net2 vss 88.1977e-18
c1370 n8__i0__i3__net2 vss 56.8403e-18
c1371 n24__rst vss 14.4474e-18
c1372 n25__rst vss 8.59666e-18
c1373 n27__rst vss 6.79178e-18
c1374 n28__rst vss 6.83761e-18
c1375 n30__rst vss 6.94772e-18
c1376 n31__rst vss 15.2238e-18
c1377 n2__net7 vss 9.84983e-18
c1378 n2__net11 vss 11.0715e-18
c1379 n30__net4 vss 17.9759e-18
c1380 n31__net4 vss 7.29803e-18
c1381 n33__net4 vss 9.08929e-18
c1382 n34__net4 vss 6.46747e-18
c1383 n36__net4 vss 7.07438e-18
c1384 n37__net4 vss 15.5257e-18
c1385 n2__i7__net5 vss 18.6627e-18
c1386 n3__i7__net5 vss 9.59616e-18
c1387 n2__i6__net5 vss 19.3232e-18
c1388 n3__i6__net5 vss 9.66976e-18
c1389 n2__i4__net5 vss 18.8947e-18
c1390 n3__i4__net5 vss 10.0184e-18
c1391 n2__i5__net5 vss 18.8324e-18
c1392 n3__i5__net5 vss 8.57272e-18
c1393 n5__x_out_b_3 vss 42.2924e-18
c1394 n5__x_out_b_2 vss 41.7567e-18
c1395 n5__x_out_b_1 vss 41.7676e-18
c1396 n5__x_out_b_0 vss 41.7567e-18
c1397 n26__i0__net1 vss 39.8962e-18
c1398 n19__i0__net8 vss 40.334e-18
c1399 n65__net10 vss 33.3343e-18
c1400 n67__net10 vss 53.8676e-18
c1401 n68__net10 vss 54.1248e-18
c1402 n71__net10 vss 33.3343e-18
c1403 n73__net10 vss 53.8676e-18
c1404 n74__net10 vss 54.1248e-18
c1405 n31__i0__net1 vss 36.4046e-18
c1406 n6__net7 vss 16.2672e-18
c1407 n7__net7 vss 6.89828e-18
c1408 n9__net7 vss 6.89965e-18
c1409 n10__net7 vss 6.93304e-18
c1410 n12__net7 vss 7.11942e-18
c1411 n13__net7 vss 16.062e-18
c1412 n6__net11 vss 17.4657e-18
c1413 n7__net11 vss 6.43843e-18
c1414 n9__net11 vss 7.16786e-18
c1415 n10__net11 vss 6.56841e-18
c1416 n12__net11 vss 8.26408e-18
c1417 n13__net11 vss 17.3916e-18
c1418 n2__y_out_b_3 vss 9.26268e-18
c1419 n2__y_out_b_2 vss 9.36511e-18
c1420 n2__y_out_b_1 vss 9.30973e-18
c1421 n2__y_out_b_0 vss 9.28398e-18
c1422 n13__i0__net9 vss 52.6078e-18
c1423 n14__i0__net9 vss 33.6404e-18
c1424 n37__net3 vss 45.6603e-18
c1425 n39__net3 vss 42.9791e-18
c1426 n41__net3 vss 44.2401e-18
c1427 n42__net3 vss 45.3844e-18
c1428 n43__net3 vss 45.6603e-18
c1429 n45__net3 vss 43.9582e-18
c1430 n47__net3 vss 43.2688e-18
c1431 n48__net3 vss 45.3844e-18
c1432 n13__i0__net10 vss 32.9673e-18
c1433 n14__i0__net10 vss 52.5306e-18
c1434 n6__i7__net2 vss 88.2839e-18
c1435 n7__i7__net2 vss 62.171e-18
c1436 n6__i6__net2 vss 88.7153e-18
c1437 n7__i6__net2 vss 62.0979e-18
c1438 n6__i4__net2 vss 88.2866e-18
c1439 n7__i4__net2 vss 62.3952e-18
c1440 n6__i5__net2 vss 88.7037e-18
c1441 n7__i5__net2 vss 61.7566e-18
c1442 n5__y_out_b_3 vss 41.8044e-18
c1443 n5__y_out_b_2 vss 42.0632e-18
c1444 n5__y_out_b_1 vss 42.0728e-18
c1445 n5__y_out_b_0 vss 41.8045e-18
c1446 n14__vdd vss 29.6871e-18
c1447 n15__vdd vss 53.0575e-18
c1448 n18__vdd vss 28.4126e-18
c1449 n19__vdd vss 36.4751e-18
c1450 n20__vdd vss 22.464e-18
c1451 n21__vdd vss 40.5729e-18
c1452 n23__vdd vss 90.7564e-18
c1453 n24__vdd vss 30.284e-18
c1454 n39__vdd vss 61.081e-18
c1455 n40__vdd vss 59.3291e-18
c1456 n46__vdd vss 48.5692e-18
c1457 n48__vdd vss 58.742e-18
c1458 n49__vdd vss 26.565e-18
c1459 n54__vdd vss 83.9784e-18
c1460 n59__vdd vss 73.0727e-18
c1461 n61__vdd vss 7.01366e-18
c1462 n64__vdd vss 28.5177e-18
c1463 n67__vdd vss 34.7087e-18
c1464 n70__vdd vss 57.6092e-18
c1465 n73__vdd vss 40.0343e-18
c1466 n76__vdd vss 63.7958e-18
c1467 n80__vdd vss 31.2383e-18
c1468 n83__vdd vss 86.445e-18
c1469 n86__vdd vss 143.649e-18
c1470 n90__vdd vss 113.925e-18
c1471 n95__vdd vss 71.1876e-18
c1472 n96__vdd vss 34.61e-18
c1473 n99__vdd vss 32.058e-18
c1474 n100__vdd vss 49.3711e-18
c1475 n101__vdd vss 39.0358e-18
c1476 n102__vdd vss 107.923e-18
c1477 n104__vdd vss 27.9856e-18
c1478 n105__vdd vss 87.5519e-18
c1479 n106__vdd vss 172.443e-18
c1480 n108__vdd vss 36.8237e-18
c1481 n109__vdd vss 36.1973e-18
c1482 n110__vdd vss 27.829e-18
c1483 n111__vdd vss 43.5367e-18
c1484 n112__vdd vss 30.3235e-18
c1485 n142__vdd vss 72.9485e-18
c1486 n145__vdd vss 54.2067e-18
c1487 n149__vdd vss 268.549e-18
c1488 n155__vdd vss 71.1864e-18
c1489 n156__vdd vss 33.7893e-18
c1490 n159__vdd vss 32.078e-18
c1491 n160__vdd vss 49.3711e-18
c1492 n161__vdd vss 38.7314e-18
c1493 n162__vdd vss 107.923e-18
c1494 n164__vdd vss 27.9682e-18
c1495 n165__vdd vss 87.5328e-18
c1496 n166__vdd vss 172.409e-18
c1497 n168__vdd vss 36.8237e-18
c1498 n169__vdd vss 36.2534e-18
c1499 n170__vdd vss 27.5556e-18
c1500 n171__vdd vss 43.5648e-18
c1501 n172__vdd vss 30.3422e-18
c1502 n202__vdd vss 72.9736e-18
c1503 n205__vdd vss 54.2704e-18
c1504 n209__vdd vss 268.601e-18
c1505 n26__i0__net8 vss 102.642e-18
c1506 n16__i0__net11 vss 98.1193e-18
c1507 n17__i0__net11 vss 141.92e-18
rd2 vdd n222__vdd 122.4e-3
rd3 vdd n220__vdd 122.4e-3
rd4 vss n252__vss 61.19e-3
rd5 n252__vss n253__vss 122.4e-3
rd6 vss n251__vss 61.19e-3
rd7 n251__vss n250__vss 122.4e-3
re1 n220__vdd n217__vdd 83.33e-3
re2 n218__vdd vdd 83.33e-3
re3 n222__vdd n219__vdd 83.33e-3
re4 n250__vss n246__vss 83.33e-3
re5 n247__vss n251__vss 83.33e-3
re6 n252__vss n248__vss 83.33e-3
re7 n249__vss n253__vss 83.33e-3
rf1 n217__vdd n214__vdd 83.33e-3
rf2 n215__vdd n218__vdd 83.33e-3
rf3 n219__vdd n216__vdd 83.33e-3
rf4 n246__vss n242__vss 83.33e-3
rf5 n243__vss n247__vss 83.33e-3
rf6 n248__vss n244__vss 83.33e-3
rf7 n245__vss n249__vss 83.33e-3
rg1 n214__vdd n10__vdd 83.33e-3
rg2 n11__vdd n215__vdd 83.33e-3
rg3 n216__vdd n12__vdd 83.33e-3
rg4 n242__vss n238__vss 83.33e-3
rg5 n239__vss n243__vss 83.33e-3
rg6 n244__vss n240__vss 83.33e-3
rg7 n241__vss n245__vss 83.33e-3
rh1 x_in_3 n5__x_in_3 40.41e-3
rh2 x_in_2 n4__x_in_2 40.41e-3
rh3 x_in_1 n5__x_in_1 40.41e-3
rh4 x_in_0 n4__x_in_0 40.41e-3
rh5 n7__vdd n10__vdd 83.33e-3
rh6 n11__vdd n8__vdd 83.33e-3
rh7 n9__vdd n12__vdd 83.33e-3
rh8 n14__i0__net7 n8__i0__net7 1.7356
rh9 n22__i0__net1 n12__i0__net1 2.6332
rh10 n23__i0__net1 n21__i0__net1 752.6e-3
rh11 n1__y_in_3 y_in_3 1.5312
rh12 n2__y_in_2 y_in_2 1.5312
rh13 n1__y_in_1 y_in_1 1.5312
rh14 n2__y_in_0 y_in_0 1.5312
rh15 n16__i0__net7 n13__i0__net7 655.2e-3
rh16 n46__rst n13__rst 3.5072
rh17 n238__vss n234__vss 83.33e-3
rh18 n235__vss n239__vss 83.33e-3
rh19 n240__vss n236__vss 83.33e-3
rh20 n237__vss n241__vss 83.33e-3
rh21 n68__net4 n10__net4 3.4562
rh22 n69__net4 n11__net4 3.4562
rh23 n70__net4 n14__net4 3.4562
rh24 n71__net4 n15__net4 3.4562
rh25 n68__net3 n64__net3 1.6055
rh26 n64__net3 n25__net3 3.3957
rh27 n69__net3 n65__net3 1.6055
rh28 n65__net3 n26__net3 3.3957
rh29 n70__net3 n66__net3 1.6055
rh30 n66__net3 n27__net3 3.3957
rh31 n71__net3 n67__net3 1.1055
rh32 n67__net3 n28__net3 3.3957
rh33 n93__net9 n89__net9 2.2851
rh34 n89__net9 n29__net9 3.2063
rh35 n94__net9 n90__net9 2.2851
rh36 n90__net9 n30__net9 3.2063
rh37 n95__net9 n91__net9 2.2851
rh38 n91__net9 n31__net9 3.2063
rh39 n96__net9 n92__net9 1.7851
rh40 n92__net9 n32__net9 3.2063
rh41 n7__x_out_3 n5__x_out_3 2.4191
rh42 n6__x_out_2 n5__x_out_2 2.4191
rh43 n7__x_out_1 n5__x_out_1 2.4191
rh44 n6__x_out_0 n5__x_out_0 2.4191
rh45 n11__x_out_b_3 n10__x_out_b_3 2.9518
rh46 n12__x_out_b_2 n9__x_out_b_2 2.9518
rh47 n11__x_out_b_1 n10__x_out_b_1 2.9518
rh48 n12__x_out_b_0 n9__x_out_b_0 2.9518
rh49 n39__net7 n38__net7 200.8e-3
rh50 n38__net7 n37__net7 712.7e-3
rh51 n38__net11 n37__net11 200.8e-3
rh52 n37__net11 n36__net11 717.6e-3
rh53 n109__net10 n105__net10 3.0616
rh54 n105__net10 n37__net10 3.0206
rh55 n110__net10 n106__net10 3.0616
rh56 n106__net10 n38__net10 3.0206
rh57 n111__net10 n107__net10 3.0616
rh58 n107__net10 n39__net10 3.0206
rh59 n112__net10 n108__net10 2.5616
rh60 n108__net10 n40__net10 3.0206
rh61 y_out_3 n5__y_out_3 61.23e-3
rh62 y_out_2 n5__y_out_2 61.23e-3
rh63 y_out_1 n5__y_out_1 61.23e-3
rh64 y_out_0 n5__y_out_0 61.23e-3
rh65 y_out_b_3 n10__y_out_b_3 136.2e-3
rh66 y_out_b_2 n10__y_out_b_2 136.2e-3
rh67 y_out_b_1 n10__y_out_b_1 136.2e-3
rh68 y_out_b_0 n10__y_out_b_0 136.2e-3
rh69 x_out_b_3 n12__x_out_b_3 308.9e-3
rh70 x_out_b_2 n11__x_out_b_2 308.9e-3
rh71 x_out_b_1 n12__x_out_b_1 308.9e-3
rh72 x_out_b_0 n11__x_out_b_0 308.9e-3
rh73 x_out_3 n6__x_out_3 344.4e-3
rh74 x_out_2 n7__x_out_2 344.4e-3
rh75 x_out_1 n6__x_out_1 344.4e-3
rh76 x_out_0 n7__x_out_0 344.4e-3
ri1 n4__x_in_3 n5__x_in_3 1
ri2 n4__x_in_2 n5__x_in_2 1
ri3 n4__x_in_1 n5__x_in_1 1
ri4 n4__x_in_0 n5__x_in_0 1
ri5 n12__rst n13__rst 1.1391
ri6 n14__rst n15__rst 1.9849
ri7 n8__i0__net6 n9__i0__net6 2.1897
ri8 n8__i0__net1 n9__i0__net1 1.2901
ri9 n4__i0__net8 n5__i0__net8 1.3196
ri11 n12__i0__net1 n13__i0__net1 500e-3
ri12 n21__net9 n29__net9 1
ri13 n30__net9 n23__net9 1
ri14 n25__net9 n31__net9 1
ri15 n32__net9 n27__net9 1
ri16 n8__i0__net7 n9__i0__net7 1
ri17 n37__net10 n29__net10 1
ri18 n31__net10 n38__net10 1
ri19 n39__net10 n33__net10 1
ri20 n35__net10 n40__net10 1
ri21 n25__net3 n21__net3 500e-3
ri22 n22__net3 n26__net3 500e-3
ri23 n27__net3 n23__net3 500e-3
ri24 n24__net3 n28__net3 500e-3
ri25 n2__vdd n7__vdd 83.33e-3
ri26 n8__vdd n3__vdd 83.33e-3
ri27 n6__vdd n9__vdd 83.33e-3
ri28 n9__net4 n10__net4 1
ri29 n11__net4 n12__net4 1
ri30 n13__net4 n14__net4 1
ri31 n15__net4 n16__net4 1
ri32 n13__i0__net7 n14__i0__net7 1.1909
ri33 n21__i0__net1 n22__i0__net1 1.3262
ri34 n9__x_out_b_3 n10__x_out_b_3 1
ri35 n9__x_out_b_2 n10__x_out_b_2 1
ri36 n9__x_out_b_1 n10__x_out_b_1 1
ri37 n9__x_out_b_0 n10__x_out_b_0 1
ri38 n4__x_out_3 n5__x_out_3 789.9e-3
ri39 n5__x_out_2 n4__x_out_2 789.9e-3
ri40 n4__x_out_1 n5__x_out_1 789.9e-3
ri41 n5__x_out_0 n4__x_out_0 789.9e-3
ri42 n18__i0__net8 n17__i0__net8 765.8e-3
ri43 n24__i0__net1 n25__i0__net1 277.8e-3
ri44 n25__i0__net1 n23__i0__net1 394.3e-3
ri45 n1__y_in_3 n2__y_in_3 1.2813
ri46 n1__y_in_2 n2__y_in_2 1.2813
ri47 n1__y_in_1 n2__y_in_1 1.2813
ri48 n1__y_in_0 n2__y_in_0 1.2813
ri49 n15__i0__net7 n16__i0__net7 1.4306
ri50 n8__i0__net11 n9__i0__net11 1.3503
ri51 n22__i0__net10 n19__i0__net10 757.2e-3
ri52 n89__net9 n62__net9 1
ri53 n64__net9 n90__net9 1
ri54 n91__net9 n66__net9 1
ri55 n68__net9 n92__net9 1
ri56 n21__i0__net9 n19__i0__net9 1.3683
ri57 n105__net10 n78__net10 1
ri58 n79__net10 n106__net10 1
ri59 n107__net10 n82__net10 1
ri60 n83__net10 n108__net10 1
ri61 n45__rst n46__rst 1.1843
ri62 n64__net3 n58__net3 500e-3
ri63 n59__net3 n65__net3 500e-3
ri64 n66__net3 n60__net3 500e-3
ri65 n61__net3 n67__net3 500e-3
ri66 n234__vss n230__vss 83.33e-3
ri67 n231__vss n235__vss 83.33e-3
ri68 n236__vss n232__vss 83.33e-3
ri69 n233__vss n237__vss 83.33e-3
ri70 n64__net4 n67__net4 775.3e-3
ri71 n67__net4 n68__net4 490.7e-3
ri73 n68__net4 n69__net4 1.0061
ri75 n69__net4 n70__net4 387.6e-3
ri77 n70__net4 n71__net4 1.0061
ri79 n36__net11 n32__net11 1.6083
ri80 n37__net7 n34__net7 500e-3
ri81 n62__net3 n68__net3 952.3e-3
ri82 n68__net3 n69__net3 861.1e-3
ri83 n69__net3 n70__net3 532.6e-3
ri84 n70__net3 n71__net3 1.3611
ri85 n86__net9 n93__net9 1.3462
ri86 n93__net9 n94__net9 721.6e-3
ri87 n94__net9 n95__net9 677.5e-3
ri88 n95__net9 n96__net9 1.2216
ri89 n6__x_out_3 n7__x_out_3 1.2115
ri90 n6__x_out_2 n7__x_out_2 1.2115
ri91 n6__x_out_1 n7__x_out_1 1.2115
ri92 n6__x_out_0 n7__x_out_0 1.2115
ri93 n11__x_out_b_3 n12__x_out_b_3 1.1363
ri94 n11__x_out_b_2 n12__x_out_b_2 1.1363
ri95 n11__x_out_b_1 n12__x_out_b_1 1.1363
ri96 n11__x_out_b_0 n12__x_out_b_0 1.1363
ri97 n35__net7 n38__net7 500e-3
ri98 n37__net11 n34__net11 500e-3
ri99 n9__y_out_b_3 n10__y_out_b_3 500e-3
ri100 n10__y_out_b_2 n9__y_out_b_2 500e-3
ri101 n9__y_out_b_1 n10__y_out_b_1 500e-3
ri102 n10__y_out_b_0 n9__y_out_b_0 500e-3
ri103 n36__net7 n39__net7 500e-3
ri104 n38__net11 n35__net11 500e-3
ri105 n4__y_out_3 n5__y_out_3 500e-3
ri106 n5__y_out_2 n4__y_out_2 500e-3
ri107 n4__y_out_1 n5__y_out_1 500e-3
ri108 n5__y_out_0 n4__y_out_0 500e-3
ri109 n102__net10 n109__net10 678.3e-3
ri110 n109__net10 n110__net10 426.3e-3
ri111 n110__net10 n111__net10 984.6e-3
ri112 n111__net10 n112__net10 926.3e-3
rj1 n4__x_in_3 n2__x_in_3 500e-3
rj2 n2__x_in_2 n5__x_in_2 500e-3
rj3 n4__x_in_1 n2__x_in_1 500e-3
rj4 n2__x_in_0 n5__x_in_0 500e-3
rj5 n9__i0__net1 n6__i0__net1 561.2e-3
rj6 n5__i0__net8 n2__i0__net8 561.2e-3
rj8 n21__net9 n17__net9 486.1e-3
rj10 n23__net9 n18__net9 486.1e-3
rj12 n25__net9 n19__net9 486.1e-3
rj14 n27__net9 n20__net9 486.1e-3
rj16 n29__net10 n18__net10 1.0759
rj18 n31__net10 n22__net10 1.0759
rj20 n33__net10 n24__net10 1.0759
rj22 n35__net10 n28__net10 1.0759
rj23 n18__i0__net1 n13__i0__net1 938.4e-3
rj24 n13__i0__net1 n10__i0__net1 47.62e-3
rj25 n9__i0__net3 n8__i0__net3 986.1e-3
rj26 n8__i0__net3 n6__i0__net3 722.8e-3
rj27 n21__net3 n10__net3 1
rj28 n12__net3 n22__net3 1
rj29 n23__net3 n16__net3 1
rj30 n18__net3 n24__net3 1
rj31 n10__i0__net7 n9__i0__net7 379.9e-3
rj32 n9__i0__net7 n7__i0__net7 695.9e-3
rj33 n16__clk clk 488.8e-3
rj34 clk n17__clk 87.08e-3
rj35 n17__clk n8__clk 830.3e-3
rj36 n13__clk n17__clk 500e-3
rj37 n16__i1__net1 n14__i1__net1 671.4e-3
rj38 n14__i1__net1 n11__i1__net1 1.1534
rj39 n16__i2__net1 n14__i2__net1 671.4e-3
rj40 n14__i2__net1 n11__i2__net1 1.1534
rj41 n16__i3__net1 n14__i3__net1 671.4e-3
rj42 n14__i3__net1 n11__i3__net1 1.1534
rj43 n16__i8__net1 n14__i8__net1 671.4e-3
rj44 n14__i8__net1 n11__i8__net1 1.1534
rj45 n17__rst n14__rst 1.6222
rj46 n19__rst rst 1.1328
rj47 rst n15__rst 484.6e-3
rj48 n15__rst rst 32.17e-3
rj49 rst n22__rst 44.08e-3
rj50 n22__rst n12__rst 4.898e-3
rj51 n8__rst n22__rst 500e-3
rj52 n5__i1__net2 n4__i1__net2 1.2984
rj53 n5__i2__net2 n4__i2__net2 1.2984
rj54 n5__i3__net2 n4__i3__net2 1.2984
rj55 n5__i8__net2 n4__i8__net2 1.2984
rj56 n16__i0__i2__net1 n14__i0__i2__net1 671.4e-3
rj57 n14__i0__i2__net1 n11__i0__i2__net1 1.1534
rj58 n16__i0__i3__net1 n14__i0__i3__net1 671.4e-3
rj59 n14__i0__i3__net1 n11__i0__i3__net1 1.1534
rj60 n5__i0__i2__net2 n4__i0__i2__net2 1.2984
rj61 n5__i0__i3__net2 n4__i0__i3__net2 1.2984
rj62 n45__net9 n41__net9 741.9e-3
rj63 n46__net9 n42__net9 741.9e-3
rj64 n47__net9 n43__net9 741.9e-3
rj65 n48__net9 n44__net9 741.9e-3
rj66 n53__net10 n49__net10 840.3e-3
rj67 n54__net10 n50__net10 840.3e-3
rj68 n55__net10 n51__net10 840.3e-3
rj69 n56__net10 n52__net10 840.3e-3
rj70 n11__i0__net3 n10__i0__net3 741.9e-3
rj71 n20__i0__net1 n19__i0__net1 741.9e-3
rj72 n18__clk n15__clk 840.3e-3
rj73 n12__i0__net7 n11__i0__net7 840.3e-3
rj74 n1__vdd n2__vdd 166.7e-3
rj75 n3__vdd n4__vdd 166.7e-3
rj76 n5__vdd n6__vdd 166.7e-3
rj77 n17__net4 n9__net4 632.8e-3
rj78 n18__net4 n12__net4 632.8e-3
rj79 n19__net4 n13__net4 632.8e-3
rj80 n20__net4 n16__net4 632.8e-3
rj81 n14__i1__net5 n11__i1__net5 1.4531
rj82 n14__i2__net5 n11__i2__net5 1.4531
rj83 n14__i3__net5 n11__i3__net5 1.4531
rj84 n14__i8__net5 n11__i8__net5 1.4531
rj85 n10__i0__net6 n8__i0__net6 2.7526
rj86 n11__i0__net6 n9__i0__net6 2.7533
rj87 n9__i0__net6 n6__i0__net6 555.8e-3
rj88 n12__i1__net4 n7__i1__net4 531.4e-3
rj89 n12__i2__net4 n7__i2__net4 531.4e-3
rj90 n12__i3__net4 n7__i3__net4 531.4e-3
rj91 n12__i8__net4 n7__i8__net4 531.4e-3
rj92 n14__i0__i2__net5 n11__i0__i2__net5 1.4531
rj93 n14__i0__i3__net5 n11__i0__i3__net5 1.4531
rj94 n13__i1__net4 n9__i1__net4 715.5e-3
rj95 n13__i2__net4 n9__i2__net4 715.5e-3
rj96 n13__i3__net4 n9__i3__net4 715.5e-3
rj97 n13__i8__net4 n9__i8__net4 715.5e-3
rj98 n12__i0__i2__net4 n7__i0__i2__net4 531.4e-3
rj99 n12__i0__i3__net4 n7__i0__i3__net4 531.4e-3
rj100 n13__i0__i2__net4 n9__i0__i2__net4 1.2155
rj101 n13__i0__i3__net4 n9__i0__i3__net4 1.2155
rj102 n17__i0__net8 n4__i0__net8 3.1053
rj103 n4__x_out_3 n2__x_out_3 1
rj104 n2__x_out_2 n4__x_out_2 1
rj105 n4__x_out_1 n2__x_out_1 1
rj106 n2__x_out_0 n4__x_out_0 1
rj107 n9__x_out_b_3 n6__x_out_b_3 617.6e-3
rj108 n10__x_out_b_2 n7__x_out_b_2 617.6e-3
rj109 n9__x_out_b_1 n6__x_out_b_1 617.6e-3
rj110 n10__x_out_b_0 n7__x_out_b_0 617.6e-3
rj111 n24__i0__net1 n8__i0__net1 3.1121
rj112 n4__y_in_3 n2__y_in_3 500e-3
rj113 n1__y_in_2 n4__y_in_2 500e-3
rj114 n4__y_in_1 n2__y_in_1 500e-3
rj115 n1__y_in_0 n4__y_in_0 500e-3
rj116 n15__i0__net7 n18__i0__net7 500e-3
rj117 n11__i0__net11 n9__i0__net11 500e-3
rj119 n31__i0__net1 n25__i0__net1 500e-3
rj120 n27__i0__net1 n31__i0__net1 500e-3
rj121 n19__i0__net10 n8__i0__net10 1
rj123 n62__net9 n57__net9 486.1e-3
rj125 n64__net9 n58__net9 486.1e-3
rj127 n66__net9 n59__net9 486.1e-3
rj129 n68__net9 n60__net9 486.1e-3
rj130 n19__i0__net9 n11__i0__net9 1
rj132 n78__net10 n66__net10 1.0759
rj134 n79__net10 n70__net10 1.0759
rj136 n82__net10 n72__net10 1.0759
rj138 n83__net10 n76__net10 1.0759
rj139 n58__net3 n38__net3 1
rj140 n40__net3 n59__net3 1
rj141 n60__net3 n44__net3 1
rj142 n46__net3 n61__net3 1
rj143 n16__i7__net1 n14__i7__net1 171.4e-3
rj144 n14__i7__net1 n11__i7__net1 1.1534
rj145 n16__i6__net1 n14__i6__net1 171.4e-3
rj146 n14__i6__net1 n11__i6__net1 1.1534
rj147 n16__i4__net1 n14__i4__net1 171.4e-3
rj148 n14__i4__net1 n11__i4__net1 1.1534
rj149 n16__i5__net1 n14__i5__net1 171.4e-3
rj150 n14__i5__net1 n11__i5__net1 1.1534
rj151 n12__i7__net2 n4__i7__net2 798.4e-3
rj152 n12__i6__net2 n4__i6__net2 798.4e-3
rj153 n12__i4__net2 n4__i4__net2 798.4e-3
rj154 n12__i5__net2 n4__i5__net2 798.4e-3
rj155 n230__vss n17__vss 166.7e-3
rj156 n63__vss n231__vss 166.7e-3
rj157 n232__vss n140__vss 166.7e-3
rj158 n198__vss n233__vss 166.7e-3
rj159 n44__rst n43__rst 204.7e-3
rj160 n43__rst n45__rst 698.9e-3
rj161 n25__i0__net8 n24__i0__net8 631.9e-3
rj162 n24__i0__net8 n26__i0__net8 237.4e-3
rj163 n26__i0__net8 n27__i0__net8 439.6e-3
rj164 n26__i0__net8 n23__i0__net8 39.63e-3
rj165 n27__i0__net8 n18__i0__net8 9.391e-3
rj166 n21__i0__net8 n27__i0__net8 500e-3
rj167 n15__i0__net11 n16__i0__net11 758.3e-3
rj168 n16__i0__net11 n17__i0__net11 602.5e-3
rj169 n17__i0__net11 n8__i0__net11 286.1e-3
rj170 n16__i0__net11 n14__i0__net11 41e-3
rj171 n17__i0__net11 n13__i0__net11 513.3e-3
rj172 n17__i0__net10 n20__i0__net10 764.3e-3
rj173 n20__i0__net10 n21__i0__net10 208.7e-3
rj174 n21__i0__net10 n22__i0__net10 956e-3
rj175 n15__i0__net10 n20__i0__net10 500e-3
rj176 n10__i0__net10 n21__i0__net10 500e-3
rj177 n17__i0__net9 n20__i0__net9 703.4e-3
rj178 n20__i0__net9 n21__i0__net9 101.9e-3
rj179 n21__i0__net9 n9__i0__net9 650.1e-3
rj180 n12__i0__net9 n20__i0__net9 500e-3
rj181 n69__net9 n61__net9 741.9e-3
rj182 n70__net9 n63__net9 741.9e-3
rj183 n71__net9 n65__net9 741.9e-3
rj184 n72__net9 n67__net9 741.9e-3
rj185 n85__net10 n77__net10 840.3e-3
rj186 n86__net10 n80__net10 840.3e-3
rj187 n87__net10 n81__net10 840.3e-3
rj188 n88__net10 n84__net10 840.3e-3
rj189 n64__net4 n65__net4 764.9e-3
rj190 n65__net4 n66__net4 197.8e-3
rj191 n66__net4 n50__net4 696.4e-3
rj192 n56__net4 n65__net4 500e-3
rj193 n53__net4 n66__net4 500e-3
rj194 n30__net7 n28__net7 923.6e-3
rj196 n29__net7 n34__net7 1
rj197 n29__net11 n32__net11 206.4e-3
rj198 n32__net11 n28__net11 1.1933
rj200 n59__net4 n58__net4 204.5e-3
rj201 n58__net4 n67__net4 587.9e-3
rj202 n56__net3 n62__net3 654.4e-3
rj203 n62__net3 n63__net3 30.42e-3
rj204 n63__net3 n50__net3 698.9e-3
rj205 n53__net3 n63__net3 500e-3
rj206 n60__net4 n68__net4 1.4279
rj207 n61__net4 n69__net4 1.4279
rj208 n62__net4 n70__net4 1.4279
rj209 n63__net4 n71__net4 1.4279
rj210 n14__i7__net5 n11__i7__net5 1.4531
rj211 n14__i6__net5 n11__i6__net5 1.4531
rj212 n14__i4__net5 n11__i4__net5 1.4531
rj213 n14__i5__net5 n11__i5__net5 1.4531
rj214 n12__i7__net4 n7__i7__net4 531.4e-3
rj215 n12__i6__net4 n7__i6__net4 531.4e-3
rj216 n12__i4__net4 n7__i4__net4 531.4e-3
rj217 n12__i5__net4 n7__i5__net4 531.4e-3
rj218 n35__net7 n31__net7 500e-3
rj219 n30__net11 n34__net11 500e-3
rj220 n13__i7__net4 n9__i7__net4 715.5e-3
rj221 n13__i6__net4 n9__i6__net4 715.5e-3
rj222 n13__i4__net4 n9__i4__net4 715.5e-3
rj223 n13__i5__net4 n9__i5__net4 715.5e-3
rj224 n36__net7 n32__net7 500e-3
rj225 n31__net11 n35__net11 500e-3
rj226 n86__net9 n87__net9 742.5e-3
rj227 n87__net9 n88__net9 203.2e-3
rj228 n88__net9 n80__net9 701e-3
rj229 n74__net9 n87__net9 500e-3
rj230 n77__net9 n88__net9 500e-3
rj231 n102__net10 n103__net10 576.3e-3
rj232 n103__net10 n104__net10 203.2e-3
rj233 n104__net10 n90__net10 701e-3
rj234 n96__net10 n103__net10 500e-3
rj235 n93__net10 n104__net10 500e-3
rj236 n2__y_out_3 n4__y_out_3 1.0955
rj237 n2__y_out_2 n4__y_out_2 1.0955
rj238 n2__y_out_1 n4__y_out_1 1.0955
rj239 n2__y_out_0 n4__y_out_0 1.0955
rj240 n9__y_out_b_3 n6__y_out_b_3 1
rj241 n7__y_out_b_2 n9__y_out_b_2 1
rj242 n9__y_out_b_1 n6__y_out_b_1 1
rj243 n7__y_out_b_0 n9__y_out_b_0 1
rj244 clk_div4_out_b n4__clk_div4_out_b 495.9e-3
rj245 clk_div4_out n4__clk_div4_out 361.2e-3
rk1 n1__x_in_3 n2__x_in_3 75.3531
rk2 n2__x_in_3 n3__x_in_3 62.2408
rk3 n1__x_in_2 n2__x_in_2 62.2408
rk4 n2__x_in_2 n3__x_in_2 75.3531
rk5 n1__x_in_1 n2__x_in_1 75.3531
rk6 n2__x_in_1 n3__x_in_1 62.2408
rk7 n1__x_in_0 n2__x_in_0 62.2408
rk8 n2__x_in_0 n3__x_in_0 75.3531
rk9 n8__clk n9__clk 4.881e-3
rk10 n10__clk n11__clk 4.881e-3
rk11 n9__clk n10__clk 12.91e-3
rk12 n2__clk n11__clk 45
rk13 n8__rst n9__rst 4.881e-3
rk14 n10__rst n11__rst 4.881e-3
rk15 n9__rst n10__rst 12.91e-3
rk16 n2__rst n11__rst 45
rk17 net9 n17__net9 509.8e-3
rk18 n18__net9 n3__net9 509.8e-3
rk19 n5__net9 n19__net9 509.8e-3
rk20 n20__net9 n7__net9 509.8e-3
rk21 n17__net10 n18__net10 3.525e-3
rk22 net10 n19__net10 3.525e-3
rk23 n17__net10 n19__net10 9.761e-3
rk24 n3__net10 n20__net10 3.525e-3
rk25 n21__net10 n22__net10 3.525e-3
rk26 n20__net10 n21__net10 9.761e-3
rk27 n23__net10 n24__net10 3.525e-3
rk28 n5__net10 n25__net10 3.525e-3
rk29 n23__net10 n25__net10 9.761e-3
rk30 n7__net10 n26__net10 3.525e-3
rk31 n27__net10 n28__net10 3.525e-3
rk32 n26__net10 n27__net10 9.761e-3
rk33 n5__i0__net3 n6__i0__net3 75.2992
rk34 n6__i0__net3 n7__i0__net3 31.3175
rk35 n5__i0__net6 n6__i0__net6 31.5214
rk36 n6__i0__net6 n7__i0__net6 75.0929
rk37 n8__i1__net1 n10__i1__net1 75.4098
rk38 n10__i1__net1 n11__i1__net1 53.73e-3
rk39 n11__i1__net1 n12__i1__net1 62.2901
rk40 n11__i1__net1 n13__i1__net1 75.4571
rk41 n9__i1__net1 n10__i1__net1 62
rk42 n8__i2__net1 n10__i2__net1 75.4127
rk43 n10__i2__net1 n11__i2__net1 53.73e-3
rk44 n11__i2__net1 n12__i2__net1 75.47
rk45 n11__i2__net1 n13__i2__net1 62.3044
rk46 n9__i2__net1 n10__i2__net1 62
rk47 n8__i3__net1 n10__i3__net1 75.4098
rk48 n10__i3__net1 n11__i3__net1 53.73e-3
rk49 n11__i3__net1 n12__i3__net1 62.2901
rk50 n11__i3__net1 n13__i3__net1 75.4571
rk51 n9__i3__net1 n10__i3__net1 62
rk52 n8__i8__net1 n10__i8__net1 75.4127
rk53 n10__i8__net1 n11__i8__net1 53.73e-3
rk54 n11__i8__net1 n12__i8__net1 75.47
rk55 n11__i8__net1 n13__i8__net1 62.3044
rk56 n9__i8__net1 n10__i8__net1 62
rk57 n5__i0__net1 n6__i0__net1 75.3629
rk58 n6__i0__net1 n7__i0__net1 62.2408
rk59 i0__net8 n2__i0__net8 62.2408
rk60 n2__i0__net8 n3__i0__net8 75.3588
rk61 i0__net3 n8__i0__net3 509.8e-3
rk62 n10__i0__net1 i0__net1 509.8e-3
rk63 i1__net2 n4__i1__net2 45.9216
rk64 i2__net2 n4__i2__net2 45.9216
rk65 i3__net2 n4__i3__net2 45.9216
rk66 i8__net2 n4__i8__net2 45.9216
rk67 n12__clk n13__clk 3.525e-3
rk68 n4__clk n14__clk 3.525e-3
rk69 n12__clk n14__clk 9.761e-3
rk70 i0__net7 n5__i0__net7 3.525e-3
rk71 n6__i0__net7 n7__i0__net7 3.525e-3
rk72 n5__i0__net7 n6__i0__net7 9.761e-3
rk73 n8__i0__i2__net1 n10__i0__i2__net1 75.4098
rk74 n10__i0__i2__net1 n11__i0__i2__net1 53.73e-3
rk75 n11__i0__i2__net1 n12__i0__i2__net1 62.2901
rk76 n11__i0__i2__net1 n13__i0__i2__net1 75.4571
rk77 n9__i0__i2__net1 n10__i0__i2__net1 62
rk78 n8__i0__i3__net1 n10__i0__i3__net1 75.4127
rk79 n10__i0__i3__net1 n11__i0__i3__net1 53.73e-3
rk80 n11__i0__i3__net1 n12__i0__i3__net1 75.47
rk81 n11__i0__i3__net1 n13__i0__i3__net1 62.3044
rk82 n9__i0__i3__net1 n10__i0__i3__net1 62
rk83 i0__i2__net2 n4__i0__i2__net2 45.9216
rk84 i0__i3__net2 n4__i0__i3__net2 45.9216
rk85 n49__net10 n29__net10 1.2186
rk86 n31__net10 n50__net10 1.2186
rk87 n51__net10 n33__net10 1.2186
rk88 n35__net10 n52__net10 1.2186
rk89 n41__net9 n21__net9 1.7598
rk90 n42__net9 n23__net9 1.7598
rk91 n43__net9 n25__net9 1.7598
rk92 n44__net9 n27__net9 1.7598
rk93 n14__i1__net1 n15__i1__net1 75.8329
rk94 n14__i2__net1 n15__i2__net1 75.8329
rk95 n14__i3__net1 n15__i3__net1 75.8329
rk96 n14__i8__net1 n15__i8__net1 75.8329
rk97 n9__net3 net3 4.364e-3
rk98 n10__net3 n11__net3 4.364e-3
rk99 n9__net3 n11__net3 24.4e-3
rk100 n12__net3 n13__net3 4.364e-3
rk101 n14__net3 n3__net3 4.364e-3
rk102 n13__net3 n14__net3 24.4e-3
rk103 n15__net3 n5__net3 4.364e-3
rk104 n16__net3 n17__net3 4.364e-3
rk105 n15__net3 n17__net3 24.4e-3
rk106 n18__net3 n19__net3 4.364e-3
rk107 n20__net3 n7__net3 4.364e-3
rk108 n19__net3 n20__net3 24.4e-3
rk109 n15__clk n16__clk 1.2186
rk110 n10__i0__net7 n11__i0__net7 1.2186
rk111 n10__i0__net3 n9__i0__net3 1.2598
rk112 n19__i0__net1 n18__i0__net1 1.2598
rk113 n4__i1__net1 n16__i1__net1 240.2e-3
rk114 n4__i2__net1 n16__i2__net1 240.2e-3
rk115 n4__i3__net1 n16__i3__net1 240.2e-3
rk116 n4__i8__net1 n16__i8__net1 240.2e-3
rk117 n14__i0__i2__net1 n15__i0__i2__net1 75.8329
rk118 n14__i0__i3__net1 n15__i0__i3__net1 75.8329
rk119 n16__rst n4__rst 4.364e-3
rk120 n17__rst n18__rst 4.364e-3
rk121 n16__rst n18__rst 24.4e-3
rk122 n19__rst n20__rst 4.364e-3
rk123 n21__rst n6__rst 4.364e-3
rk124 n20__rst n21__rst 24.4e-3
rk125 n4__i0__i2__net1 n16__i0__i2__net1 240.2e-3
rk126 n4__i0__i3__net1 n16__i0__i3__net1 240.2e-3
rk127 n6__i1__net2 n7__i1__net2 75.167
rk128 n7__i1__net2 n8__i1__net2 299.2e-3
rk129 n8__i1__net2 n10__i1__net2 329.8e-3
rk130 n7__i1__net2 n11__i1__net2 62.4611
rk131 n8__i1__net2 n12__i1__net2 37.7267
rk132 n10__i1__net2 n5__i1__net2 115.7e-3
rk133 n9__i1__net2 n10__i1__net2 15.5
rk134 n6__i2__net2 n7__i2__net2 62.4611
rk135 n7__i2__net2 n8__i2__net2 299.2e-3
rk136 n8__i2__net2 n9__i2__net2 37.7267
rk137 n7__i2__net2 n10__i2__net2 75.167
rk138 n8__i2__net2 n12__i2__net2 329.8e-3
rk139 n12__i2__net2 n5__i2__net2 119.8e-3
rk140 n11__i2__net2 n12__i2__net2 15.5
rk141 n6__i3__net2 n7__i3__net2 75.167
rk142 n7__i3__net2 n8__i3__net2 299.2e-3
rk143 n8__i3__net2 n10__i3__net2 329.8e-3
rk144 n7__i3__net2 n11__i3__net2 62.4611
rk145 n8__i3__net2 n12__i3__net2 37.7267
rk146 n10__i3__net2 n5__i3__net2 115.7e-3
rk147 n9__i3__net2 n10__i3__net2 15.5
rk148 n6__i8__net2 n7__i8__net2 62.4611
rk149 n7__i8__net2 n8__i8__net2 299.2e-3
rk150 n8__i8__net2 n9__i8__net2 37.7267
rk151 n7__i8__net2 n10__i8__net2 75.167
rk152 n8__i8__net2 n12__i8__net2 329.8e-3
rk153 n12__i8__net2 n5__i8__net2 119.8e-3
rk154 n11__i8__net2 n12__i8__net2 15.5
rk155 n9__net10 n53__net10 509.8e-3
rk156 n9__net9 n45__net9 509.8e-3
rk157 n46__net9 n11__net9 509.8e-3
rk158 n54__net10 n11__net10 509.8e-3
rk159 n13__net10 n55__net10 509.8e-3
rk160 n13__net9 n47__net9 509.8e-3
rk161 n48__net9 n15__net9 509.8e-3
rk162 n56__net10 n15__net10 509.8e-3
rk163 n8__i1__net5 n10__i1__net5 75.4098
rk164 n10__i1__net5 n11__i1__net5 53.73e-3
rk165 n11__i1__net5 n12__i1__net5 62.2865
rk166 n11__i1__net5 n13__i1__net5 75.4571
rk167 n9__i1__net5 n10__i1__net5 62
rk168 n8__i2__net5 n10__i2__net5 75.4127
rk169 n10__i2__net5 n11__i2__net5 53.73e-3
rk170 n11__i2__net5 n12__i2__net5 75.47
rk171 n11__i2__net5 n13__i2__net5 62.3006
rk172 n9__i2__net5 n10__i2__net5 62
rk173 n8__i3__net5 n10__i3__net5 75.4098
rk174 n10__i3__net5 n11__i3__net5 53.73e-3
rk175 n11__i3__net5 n12__i3__net5 62.2865
rk176 n11__i3__net5 n13__i3__net5 75.4571
rk177 n9__i3__net5 n10__i3__net5 62
rk178 n8__i8__net5 n10__i8__net5 75.4127
rk179 n10__i8__net5 n11__i8__net5 53.73e-3
rk180 n11__i8__net5 n12__i8__net5 75.47
rk181 n11__i8__net5 n13__i8__net5 62.3006
rk182 n9__i8__net5 n10__i8__net5 62
rk183 n6__i0__i2__net2 n7__i0__i2__net2 75.167
rk184 n7__i0__i2__net2 n8__i0__i2__net2 299.2e-3
rk185 n8__i0__i2__net2 n10__i0__i2__net2 329.8e-3
rk186 n7__i0__i2__net2 n11__i0__i2__net2 62.4611
rk187 n8__i0__i2__net2 n12__i0__i2__net2 37.7267
rk188 n10__i0__i2__net2 n5__i0__i2__net2 115.7e-3
rk189 n9__i0__i2__net2 n10__i0__i2__net2 15.5
rk190 n6__i0__i3__net2 n7__i0__i3__net2 62.4611
rk191 n7__i0__i3__net2 n8__i0__i3__net2 299.2e-3
rk192 n8__i0__i3__net2 n9__i0__i3__net2 37.7267
rk193 n7__i0__i3__net2 n10__i0__i3__net2 75.167
rk194 n8__i0__i3__net2 n12__i0__i3__net2 329.8e-3
rk195 n12__i0__i3__net2 n5__i0__i3__net2 119.8e-3
rk196 n11__i0__i3__net2 n12__i0__i3__net2 15.5
rk197 n6__clk n18__clk 509.8e-3
rk198 n3__i0__net3 n11__i0__net3 509.8e-3
rk199 n20__i0__net1 n3__i0__net1 509.8e-3
rk200 n12__i0__net7 n3__i0__net7 509.8e-3
rk201 i1__net4 n7__i1__net4 45.9216
rk202 i2__net4 n7__i2__net4 45.9216
rk203 i3__net4 n7__i3__net4 45.9216
rk204 i8__net4 n7__i8__net4 45.9216
rk205 n8__i0__i2__net5 n10__i0__i2__net5 75.4098
rk206 n10__i0__i2__net5 n11__i0__i2__net5 53.73e-3
rk207 n11__i0__i2__net5 n12__i0__i2__net5 62.2865
rk208 n11__i0__i2__net5 n13__i0__i2__net5 75.4571
rk209 n9__i0__i2__net5 n10__i0__i2__net5 62
rk210 n8__i0__i3__net5 n10__i0__i3__net5 75.4127
rk211 n10__i0__i3__net5 n11__i0__i3__net5 53.73e-3
rk212 n11__i0__i3__net5 n12__i0__i3__net5 75.47
rk213 n11__i0__i3__net5 n13__i0__i3__net5 62.3006
rk214 n9__i0__i3__net5 n10__i0__i3__net5 62
rk215 i0__i2__net4 n7__i0__i2__net4 45.9216
rk216 i0__i3__net4 n7__i0__i3__net4 45.9216
rk217 n2__net4 n17__net4 41.38e-3
rk218 n4__net4 n18__net4 41.38e-3
rk219 n6__net4 n19__net4 41.38e-3
rk220 n8__net4 n20__net4 41.38e-3
rk221 n4__i1__net5 n14__i1__net5 221e-3
rk222 n14__i1__net5 n15__i1__net5 62.0171
rk223 n4__i2__net5 n14__i2__net5 221e-3
rk224 n14__i2__net5 n15__i2__net5 62.0171
rk225 n4__i3__net5 n14__i3__net5 221e-3
rk226 n14__i3__net5 n15__i3__net5 62.0171
rk227 n4__i8__net5 n14__i8__net5 221e-3
rk228 n14__i8__net5 n15__i8__net5 62.0171
rk229 n2__i0__net6 n10__i0__net6 41.38e-3
rk230 n4__i0__net6 n11__i0__net6 41.38e-3
rk231 n8__i1__net4 n9__i1__net4 37.7068
rk232 n9__i1__net4 n11__i1__net4 309.9e-3
rk233 n11__i1__net4 n12__i1__net4 615.7e-3
rk234 n10__i1__net4 n11__i1__net4 15.5
rk235 n8__i2__net4 n9__i2__net4 37.7068
rk236 n9__i2__net4 n11__i2__net4 309.9e-3
rk237 n11__i2__net4 n12__i2__net4 619.8e-3
rk238 n10__i2__net4 n11__i2__net4 15.5
rk239 n8__i3__net4 n9__i3__net4 37.7068
rk240 n9__i3__net4 n11__i3__net4 309.9e-3
rk241 n11__i3__net4 n12__i3__net4 615.7e-3
rk242 n10__i3__net4 n11__i3__net4 15.5
rk243 n8__i8__net4 n9__i8__net4 37.7068
rk244 n9__i8__net4 n11__i8__net4 309.9e-3
rk245 n11__i8__net4 n12__i8__net4 619.8e-3
rk246 n10__i8__net4 n11__i8__net4 15.5
rk247 n4__i0__i2__net5 n14__i0__i2__net5 221e-3
rk248 n14__i0__i2__net5 n15__i0__i2__net5 62.0171
rk249 n4__i0__i3__net5 n14__i0__i3__net5 221e-3
rk250 n14__i0__i3__net5 n15__i0__i3__net5 62.0171
rk251 n5__i1__net4 n13__i1__net4 45.5279
rk252 n5__i2__net4 n13__i2__net4 45.5279
rk253 n5__i3__net4 n13__i3__net4 45.5279
rk254 n5__i8__net4 n13__i8__net4 45.5279
rk255 n8__i0__i2__net4 n9__i0__i2__net4 37.7068
rk256 n9__i0__i2__net4 n11__i0__i2__net4 309.9e-3
rk257 n11__i0__i2__net4 n12__i0__i2__net4 615.7e-3
rk258 n10__i0__i2__net4 n11__i0__i2__net4 15.5
rk259 n8__i0__i3__net4 n9__i0__i3__net4 37.7068
rk260 n9__i0__i3__net4 n11__i0__i3__net4 309.9e-3
rk261 n11__i0__i3__net4 n12__i0__i3__net4 619.8e-3
rk262 n10__i0__i3__net4 n11__i0__i3__net4 15.5
rk263 n3__x_out_b_3 n5__x_out_b_3 124.6e-3
rk264 n5__x_out_b_3 n6__x_out_b_3 188.9e-3
rk265 n6__x_out_b_3 n7__x_out_b_3 15.6036
rk266 n5__x_out_b_3 n8__x_out_b_3 37.7229
rk267 n3__x_out_b_2 n5__x_out_b_2 124.6e-3
rk268 n5__x_out_b_2 n6__x_out_b_2 37.7229
rk269 n5__x_out_b_2 n7__x_out_b_2 188.9e-3
rk270 n7__x_out_b_2 n8__x_out_b_2 15.6036
rk271 n3__x_out_b_1 n5__x_out_b_1 124.6e-3
rk272 n5__x_out_b_1 n6__x_out_b_1 188.9e-3
rk273 n6__x_out_b_1 n7__x_out_b_1 15.6036
rk274 n5__x_out_b_1 n8__x_out_b_1 37.7229
rk275 n3__x_out_b_0 n5__x_out_b_0 124.6e-3
rk276 n5__x_out_b_0 n6__x_out_b_0 37.7229
rk277 n5__x_out_b_0 n7__x_out_b_0 188.9e-3
rk278 n7__x_out_b_0 n8__x_out_b_0 15.6036
rk279 n5__i0__i2__net4 n13__i0__i2__net4 45.0279
rk280 n5__i0__i3__net4 n13__i0__i3__net4 45.0279
rk281 n1__x_out_3 n2__x_out_3 37.6651
rk282 n2__x_out_3 n3__x_out_3 15.8309
rk283 n1__x_out_2 n2__x_out_2 15.8309
rk284 n2__x_out_2 n3__x_out_2 37.6651
rk285 n1__x_out_1 n2__x_out_1 37.6651
rk286 n2__x_out_1 n3__x_out_1 15.8309
rk287 n1__x_out_0 n2__x_out_0 15.8309
rk288 n2__x_out_0 n3__x_out_0 37.6651
rk289 n16__i0__net1 n26__i0__net1 124.6e-3
rk290 n26__i0__net1 n27__i0__net1 188.9e-3
rk291 n27__i0__net1 n28__i0__net1 15.6036
rk292 n26__i0__net1 n29__i0__net1 37.7229
rk293 n8__i0__net8 n19__i0__net8 124.6e-3
rk294 n19__i0__net8 n20__i0__net8 37.7229
rk295 n19__i0__net8 n21__i0__net8 188.9e-3
rk296 n21__i0__net8 n22__i0__net8 15.6036
rk297 n3__y_in_3 n4__y_in_3 75.3531
rk298 n4__y_in_3 n5__y_in_3 62.2408
rk299 n3__y_in_2 n4__y_in_2 62.2408
rk300 n4__y_in_2 n5__y_in_2 75.3531
rk301 n3__y_in_1 n4__y_in_1 75.3531
rk302 n4__y_in_1 n5__y_in_1 62.2408
rk303 n3__y_in_0 n4__y_in_0 62.2408
rk304 n4__y_in_0 n5__y_in_0 75.3531
rk305 n33__net9 n57__net9 509.8e-3
rk306 n58__net9 n35__net9 509.8e-3
rk307 n37__net9 n59__net9 509.8e-3
rk308 n60__net9 n39__net9 509.8e-3
rk309 n17__i0__net7 n18__i0__net7 37.6651
rk310 n18__i0__net7 n19__i0__net7 15.8309
rk311 n10__i0__net11 n11__i0__net11 15.8309
rk312 n11__i0__net11 n12__i0__net11 37.6651
rk313 n65__net10 n66__net10 3.525e-3
rk314 n41__net10 n67__net10 3.525e-3
rk315 n65__net10 n67__net10 9.761e-3
rk316 n43__net10 n68__net10 3.525e-3
rk317 n69__net10 n70__net10 3.525e-3
rk318 n68__net10 n69__net10 9.761e-3
rk319 n71__net10 n72__net10 3.525e-3
rk320 n45__net10 n73__net10 3.525e-3
rk321 n71__net10 n73__net10 9.761e-3
rk322 n47__net10 n74__net10 3.525e-3
rk323 n75__net10 n76__net10 3.525e-3
rk324 n74__net10 n75__net10 9.761e-3
rk325 n8__i7__net1 n10__i7__net1 75.4098
rk326 n10__i7__net1 n11__i7__net1 53.73e-3
rk327 n11__i7__net1 n12__i7__net1 62.2901
rk328 n11__i7__net1 n13__i7__net1 75.4571
rk329 n9__i7__net1 n10__i7__net1 62
rk330 n8__i6__net1 n10__i6__net1 75.4127
rk331 n10__i6__net1 n11__i6__net1 53.73e-3
rk332 n11__i6__net1 n12__i6__net1 75.47
rk333 n11__i6__net1 n13__i6__net1 62.3044
rk334 n9__i6__net1 n10__i6__net1 62
rk335 n8__i4__net1 n10__i4__net1 75.4098
rk336 n10__i4__net1 n11__i4__net1 53.73e-3
rk337 n11__i4__net1 n12__i4__net1 62.2901
rk338 n11__i4__net1 n13__i4__net1 75.4571
rk339 n9__i4__net1 n10__i4__net1 62
rk340 n8__i5__net1 n10__i5__net1 75.4127
rk341 n10__i5__net1 n11__i5__net1 53.73e-3
rk342 n11__i5__net1 n12__i5__net1 75.47
rk343 n11__i5__net1 n13__i5__net1 62.3044
rk344 n9__i5__net1 n10__i5__net1 62
rk345 n3__i0__net10 n8__i0__net10 1.762e-3
rk346 n11__i0__net8 n23__i0__net8 505.8e-3
rk347 i7__net2 n4__i7__net2 45.9216
rk348 i6__net2 n4__i6__net2 45.9216
rk349 i4__net2 n4__i4__net2 45.9216
rk350 i5__net2 n4__i5__net2 45.9216
rk351 n25__net11 n27__net11 38.0228
rk352 n27__net11 n28__net11 593.2e-3
rk353 n26__net11 n27__net11 15.5
rk354 n8__i0__net9 n9__i0__net9 31.3477
rk355 n9__i0__net9 n10__i0__net9 75.1026
rk356 n13__i0__net11 i0__net11 4.881e-3
rk357 n24__i0__net8 n12__i0__net8 1.4204
rk358 n3__i0__net9 n11__i0__net9 1.762e-3
rk359 n25__net7 n27__net7 16.0181
rk360 n27__net7 n28__net7 506.1e-3
rk361 n26__net7 n27__net7 37.5
rk362 n77__net10 n78__net10 1.2186
rk363 n79__net10 n80__net10 1.2186
rk364 n81__net10 n82__net10 1.2186
rk365 n83__net10 n84__net10 1.2186
rk366 n12__i0__net9 n13__i0__net9 3.99e-3
rk367 n14__i0__net9 n15__i0__net9 3.99e-3
rk368 n13__i0__net9 n14__i0__net9 17.08e-3
rk369 n6__i0__net9 n15__i0__net9 45
rk370 n61__net9 n62__net9 1.7598
rk371 n63__net9 n64__net9 1.7598
rk372 n65__net9 n66__net9 1.7598
rk373 n67__net9 n68__net9 1.7598
rk374 n9__i0__net10 n10__i0__net10 15.7236
rk375 n10__i0__net10 n11__i0__net10 37.7792
rk376 n14__i7__net1 n15__i7__net1 75.8329
rk377 n14__i6__net1 n15__i6__net1 75.8329
rk378 n14__i4__net1 n15__i4__net1 75.8329
rk379 n14__i5__net1 n15__i5__net1 75.8329
rk380 n16__i0__net9 n17__i0__net9 15.8709
rk381 n17__i0__net9 n18__i0__net9 37.6319
rk382 n49__net4 n50__net4 37.8736
rk383 n50__net4 n51__net4 15.6404
rk384 n37__net3 n29__net3 4.364e-3
rk385 n38__net3 n39__net3 4.364e-3
rk386 n37__net3 n39__net3 24.4e-3
rk387 n40__net3 n41__net3 4.364e-3
rk388 n42__net3 n31__net3 4.364e-3
rk389 n41__net3 n42__net3 24.4e-3
rk390 n43__net3 n33__net3 4.364e-3
rk391 n44__net3 n45__net3 4.364e-3
rk392 n43__net3 n45__net3 24.4e-3
rk393 n46__net3 n47__net3 4.364e-3
rk394 n48__net3 n35__net3 4.364e-3
rk395 n47__net3 n48__net3 24.4e-3
rk396 n12__i0__net10 n13__i0__net10 3.99e-3
rk397 n14__i0__net10 n15__i0__net10 3.99e-3
rk398 n13__i0__net10 n14__i0__net10 17.08e-3
rk399 n6__i0__net10 n12__i0__net10 45
rk400 n29__rst n43__rst 45.5
rk401 n4__i7__net1 n16__i7__net1 740.2e-3
rk402 n4__i6__net1 n16__i6__net1 740.2e-3
rk403 n4__i4__net1 n16__i4__net1 740.2e-3
rk404 n4__i5__net1 n16__i5__net1 740.2e-3
rk405 n52__net4 n53__net4 37.8889
rk406 n53__net4 n54__net4 15.6404
rk407 n5__i0__net11 n14__i0__net11 1.5681
rk408 n44__rst n26__rst 45.5018
rk409 n25__i0__net8 n16__i0__net8 501.9e-3
rk410 n16__i0__net10 n17__i0__net10 31.1929
rk411 n17__i0__net10 n18__i0__net10 75.2574
rk412 n55__net4 n56__net4 37.8736
rk413 n56__net4 n57__net4 15.6404
rk414 n7__i0__net11 n15__i0__net11 5.821e-3
rk415 n5__i7__net2 n6__i7__net2 75.167
rk416 n6__i7__net2 n7__i7__net2 293.4e-3
rk417 n7__i7__net2 n9__i7__net2 329.8e-3
rk418 n6__i7__net2 n10__i7__net2 62.4611
rk419 n7__i7__net2 n11__i7__net2 37.7267
rk420 n9__i7__net2 n12__i7__net2 615.7e-3
rk421 n8__i7__net2 n9__i7__net2 15.5
rk422 n5__i6__net2 n6__i6__net2 62.4611
rk423 n6__i6__net2 n7__i6__net2 299.2e-3
rk424 n7__i6__net2 n8__i6__net2 37.7267
rk425 n6__i6__net2 n9__i6__net2 75.167
rk426 n7__i6__net2 n11__i6__net2 329.8e-3
rk427 n11__i6__net2 n12__i6__net2 619.8e-3
rk428 n10__i6__net2 n11__i6__net2 15.5
rk429 n5__i4__net2 n6__i4__net2 75.167
rk430 n6__i4__net2 n7__i4__net2 299.2e-3
rk431 n7__i4__net2 n9__i4__net2 329.8e-3
rk432 n6__i4__net2 n10__i4__net2 62.4611
rk433 n7__i4__net2 n11__i4__net2 37.7267
rk434 n9__i4__net2 n12__i4__net2 615.7e-3
rk435 n8__i4__net2 n9__i4__net2 15.5
rk436 n5__i5__net2 n6__i5__net2 62.4611
rk437 n6__i5__net2 n7__i5__net2 299.2e-3
rk438 n7__i5__net2 n8__i5__net2 37.7267
rk439 n6__i5__net2 n9__i5__net2 75.167
rk440 n7__i5__net2 n11__i5__net2 329.8e-3
rk441 n11__i5__net2 n12__i5__net2 619.8e-3
rk442 n10__i5__net2 n11__i5__net2 15.5
rk443 n57__net10 n85__net10 509.8e-3
rk444 n49__net9 n69__net9 509.8e-3
rk445 n70__net9 n51__net9 509.8e-3
rk446 n86__net10 n59__net10 509.8e-3
rk447 n61__net10 n87__net10 509.8e-3
rk448 n53__net9 n71__net9 509.8e-3
rk449 n72__net9 n55__net9 509.8e-3
rk450 n88__net10 n63__net10 509.8e-3
rk451 n49__net3 n50__net3 15.9451
rk452 n50__net3 n51__net3 37.5
rk453 n8__i7__net5 n10__i7__net5 75.4098
rk454 n10__i7__net5 n11__i7__net5 53.73e-3
rk455 n11__i7__net5 n12__i7__net5 62.2865
rk456 n11__i7__net5 n13__i7__net5 75.4571
rk457 n9__i7__net5 n10__i7__net5 62
rk458 n8__i6__net5 n10__i6__net5 75.4127
rk459 n10__i6__net5 n11__i6__net5 53.73e-3
rk460 n11__i6__net5 n12__i6__net5 75.47
rk461 n11__i6__net5 n13__i6__net5 62.3006
rk462 n9__i6__net5 n10__i6__net5 62
rk463 n8__i4__net5 n10__i4__net5 75.4098
rk464 n10__i4__net5 n11__i4__net5 53.73e-3
rk465 n11__i4__net5 n12__i4__net5 62.2865
rk466 n11__i4__net5 n13__i4__net5 75.4571
rk467 n9__i4__net5 n10__i4__net5 62
rk468 n8__i5__net5 n10__i5__net5 75.4127
rk469 n10__i5__net5 n11__i5__net5 53.73e-3
rk470 n11__i5__net5 n12__i5__net5 75.47
rk471 n11__i5__net5 n13__i5__net5 62.3006
rk472 n9__i5__net5 n10__i5__net5 62
rk473 n58__net4 n35__net4 45.5018
rk474 n3__net7 n29__net7 27.92e-3
rk475 n29__net7 n30__net7 680.7e-3
rk476 i7__net4 n7__i7__net4 45.9216
rk477 i6__net4 n7__i6__net4 45.9216
rk478 i4__net4 n7__i4__net4 45.9216
rk479 i5__net4 n7__i5__net4 45.9216
rk480 n52__net3 n53__net3 15.9604
rk481 n53__net3 n54__net3 37.5
rk482 n1__clk_div4_out_b n3__clk_div4_out_b 16.0496
rk483 n3__clk_div4_out_b n4__clk_div4_out_b 504.9e-3
rk484 n2__clk_div4_out_b n3__clk_div4_out_b 37.5
rk485 n32__net4 n59__net4 45.5
rk486 n55__net3 n56__net3 15.9451
rk487 n56__net3 n57__net3 37.5
rk488 n22__net4 n60__net4 41.38e-3
rk489 n24__net4 n61__net4 41.38e-3
rk490 n26__net4 n62__net4 41.38e-3
rk491 n28__net4 n63__net4 41.38e-3
rk492 n3__net11 n29__net11 892.1e-3
rk493 n1__clk_div4_out n3__clk_div4_out 38.0044
rk494 n3__clk_div4_out n4__clk_div4_out 588.3e-3
rk495 n2__clk_div4_out n3__clk_div4_out 15.5
rk496 n4__i7__net5 n14__i7__net5 221e-3
rk497 n14__i7__net5 n15__i7__net5 62.0171
rk498 n4__i6__net5 n14__i6__net5 221e-3
rk499 n14__i6__net5 n15__i6__net5 62.0171
rk500 n4__i4__net5 n14__i4__net5 221e-3
rk501 n14__i4__net5 n15__i4__net5 62.0171
rk502 n4__i5__net5 n14__i5__net5 221e-3
rk503 n14__i5__net5 n15__i5__net5 62.0171
rk504 n8__i7__net4 n9__i7__net4 37.7068
rk505 n9__i7__net4 n11__i7__net4 309.9e-3
rk506 n11__i7__net4 n12__i7__net4 615.7e-3
rk507 n10__i7__net4 n11__i7__net4 15.5
rk508 n8__i6__net4 n9__i6__net4 37.7068
rk509 n9__i6__net4 n11__i6__net4 309.9e-3
rk510 n11__i6__net4 n12__i6__net4 619.8e-3
rk511 n10__i6__net4 n11__i6__net4 15.5
rk512 n8__i4__net4 n9__i4__net4 37.7068
rk513 n9__i4__net4 n11__i4__net4 309.9e-3
rk514 n11__i4__net4 n12__i4__net4 615.7e-3
rk515 n10__i4__net4 n11__i4__net4 15.5
rk516 n8__i5__net4 n9__i5__net4 37.7068
rk517 n9__i5__net4 n11__i5__net4 309.9e-3
rk518 n11__i5__net4 n12__i5__net4 619.8e-3
rk519 n10__i5__net4 n11__i5__net4 15.5
rk520 n73__net9 n74__net9 37.8701
rk521 n74__net9 n75__net9 15.6447
rk522 n89__net10 n90__net10 15.9451
rk523 n90__net10 n91__net10 37.5
rk524 n11__net7 n31__net7 45.5
rk525 n11__net11 n30__net11 45.5
rk526 n76__net9 n77__net9 37.8854
rk527 n77__net9 n78__net9 15.6447
rk528 n92__net10 n93__net10 15.9604
rk529 n93__net10 n94__net10 37.5
rk530 n5__i7__net4 n13__i7__net4 45.5279
rk531 n5__i6__net4 n13__i6__net4 45.5279
rk532 n5__i4__net4 n13__i4__net4 45.5279
rk533 n5__i5__net4 n13__i5__net4 45.5279
rk534 n8__net7 n32__net7 45.5
rk535 n8__net11 n31__net11 45.5
rk536 n79__net9 n80__net9 37.8701
rk537 n80__net9 n81__net9 15.6447
rk538 n95__net10 n96__net10 15.9451
rk539 n96__net10 n97__net10 37.5
rk540 n3__y_out_b_3 n5__y_out_b_3 124.6e-3
rk541 n5__y_out_b_3 n6__y_out_b_3 188.9e-3
rk542 n6__y_out_b_3 n7__y_out_b_3 15.6036
rk543 n5__y_out_b_3 n8__y_out_b_3 37.7229
rk544 n3__y_out_b_2 n5__y_out_b_2 124.6e-3
rk545 n5__y_out_b_2 n6__y_out_b_2 37.7229
rk546 n5__y_out_b_2 n7__y_out_b_2 188.9e-3
rk547 n7__y_out_b_2 n8__y_out_b_2 15.6036
rk548 n3__y_out_b_1 n5__y_out_b_1 124.6e-3
rk549 n5__y_out_b_1 n6__y_out_b_1 188.9e-3
rk550 n6__y_out_b_1 n7__y_out_b_1 15.6036
rk551 n5__y_out_b_1 n8__y_out_b_1 37.7229
rk552 n3__y_out_b_0 n5__y_out_b_0 124.6e-3
rk553 n5__y_out_b_0 n6__y_out_b_0 37.7229
rk554 n5__y_out_b_0 n7__y_out_b_0 188.9e-3
rk555 n7__y_out_b_0 n8__y_out_b_0 15.6036
rk556 n1__y_out_3 n2__y_out_3 37.6651
rk557 n2__y_out_3 n3__y_out_3 15.8309
rk558 n1__y_out_2 n2__y_out_2 15.8309
rk559 n2__y_out_2 n3__y_out_2 37.6651
rk560 n1__y_out_1 n2__y_out_1 37.6651
rk561 n2__y_out_1 n3__y_out_1 15.8309
rk562 n1__y_out_0 n2__y_out_0 15.8309
rk563 n2__y_out_0 n3__y_out_0 37.6651
rk564 n1__vss n2__vss 37.7885
rk565 n2__vss n4__vss 101.6e-3
rk566 n4__vss n5__vss 101.6e-3
rk567 n5__vss n6__vss 115e-3
rk568 n6__vss n7__vss 137.4e-3
rk569 n7__vss n8__vss 151.2e-3
rk570 n2__vss n9__vss 37.6968
rk571 n4__vss n10__vss 37.6926
rk572 n5__vss n11__vss 37.6853
rk573 n6__vss n12__vss 37.6853
rk574 n7__vss n13__vss 37.6962
rk575 n8__vss n14__vss 37.6811
rk576 n8__vss n15__vss 91.65e-3
rk577 n15__vss n16__vss 37.6968
rk578 n15__vss n17__vss 53.17e-3
rk579 n17__vss n18__vss 37.6926
rk580 n17__vss n19__vss 150e-3
rk581 n19__vss n20__vss 37.6876
rk582 n19__vss n21__vss 115e-3
rk583 n21__vss n22__vss 37.6853
rk584 n21__vss n23__vss 115e-3
rk585 n23__vss n24__vss 37.6853
rk586 n23__vss n25__vss 69.31e-3
rk587 n25__vss n26__vss 55.65e-3
rk588 n26__vss n27__vss 37.6853
rk589 n26__vss vss 30.82e-3
rk590 vss n28__vss 84.2e-3
rk591 n28__vss n29__vss 37.6853
rk592 n28__vss n30__vss 64.12e-3
rk593 n30__vss n31__vss 37.6853
rk594 n30__vss n32__vss 101.4e-3
rk595 n32__vss n33__vss 37.6853
rk596 n32__vss n34__vss 82.74e-3
rk597 n34__vss n35__vss 75.2174
rk598 n34__vss n36__vss 174.8e-3
rk599 n36__vss n37__vss 186e-3
rk600 n37__vss n38__vss 37.6853
rk601 n37__vss n39__vss 101.4e-3
rk602 n39__vss n40__vss 37.6853
rk603 n39__vss n41__vss 64.12e-3
rk604 n41__vss n42__vss 75.222
rk605 n41__vss n43__vss 115e-3
rk606 n43__vss n44__vss 75.2196
rk607 n43__vss n45__vss 127.7e-3
rk608 n45__vss n46__vss 75.4156
rk609 n3__vss n4__vss 4.4286
rk610 n3__vss n8__vss 3.1
rk611 n3__vss n25__vss 3.1
rk612 n3__vss n36__vss 3.1
rk613 n3__vss n45__vss 3.1
rk614 n13__vdd n14__vdd 15.8447
rk615 n14__vdd n15__vdd 94.04e-3
rk616 n15__vdd n17__vdd 101.4e-3
rk617 n17__vdd n18__vdd 101.4e-3
rk618 n18__vdd n19__vdd 58.93e-3
rk619 n19__vdd n20__vdd 55.43e-3
rk620 n20__vdd n21__vdd 45.49e-3
rk621 n21__vdd n22__vdd 89.07e-3
rk622 n22__vdd n23__vdd 12.09e-3
rk623 n23__vdd n24__vdd 101.4e-3
rk624 n24__vdd n25__vdd 39.51e-3
rk625 n14__vdd n26__vdd 15.8188
rk626 n15__vdd n27__vdd 15.8926
rk627 n15__vdd n28__vdd 15.8926
rk628 n17__vdd n29__vdd 15.7958
rk629 n17__vdd n30__vdd 15.7958
rk630 n18__vdd n31__vdd 15.8791
rk631 n18__vdd n32__vdd 15.8773
rk632 n19__vdd n33__vdd 15.7864
rk633 n20__vdd n34__vdd 15.7933
rk634 n21__vdd n35__vdd 15.8
rk635 n22__vdd n36__vdd 15.786
rk636 n23__vdd n37__vdd 15.8
rk637 n24__vdd n38__vdd 15.777
rk638 n25__vdd n39__vdd 91.65e-3
rk639 n39__vdd n40__vdd 36.8e-3
rk640 n40__vdd n42__vdd 421.3e-3
rk641 n42__vdd n43__vdd 75.5355
rk642 n25__vdd n44__vdd 15.7728
rk643 n39__vdd n45__vdd 15.8
rk644 n40__vdd n46__vdd 63.9e-3
rk645 n46__vdd n47__vdd 15.9086
rk646 n46__vdd n48__vdd 101.1e-3
rk647 n48__vdd n49__vdd 64.12e-3
rk648 n49__vdd n50__vdd 15.7967
rk649 n46__vdd n51__vdd 15.8926
rk650 n48__vdd n52__vdd 15.777
rk651 n49__vdd n53__vdd 49.87e-3
rk652 n53__vdd n54__vdd 13.87e-3
rk653 n54__vdd n56__vdd 380e-3
rk654 n56__vdd n57__vdd 75.5355
rk655 n53__vdd n58__vdd 15.782
rk656 n54__vdd n59__vdd 101.4e-3
rk657 n59__vdd n60__vdd 69.31e-3
rk658 n60__vdd n61__vdd 55.43e-3
rk659 n61__vdd n62__vdd 15.8697
rk660 n59__vdd n63__vdd 15.777
rk661 n61__vdd vdd 30.6e-3
rk662 vdd n64__vdd 83.99e-3
rk663 n64__vdd n65__vdd 15.8697
rk664 n61__vdd n66__vdd 15.8697
rk665 n64__vdd n67__vdd 63.68e-3
rk666 n67__vdd n68__vdd 15.8697
rk667 n64__vdd n69__vdd 15.8697
rk668 n67__vdd n70__vdd 100.9e-3
rk669 n70__vdd n71__vdd 15.8697
rk670 n67__vdd n72__vdd 15.8697
rk671 n70__vdd n73__vdd 114.6e-3
rk672 n73__vdd n74__vdd 62.4805
rk673 n70__vdd n75__vdd 15.8697
rk674 n73__vdd n76__vdd 63.68e-3
rk675 n76__vdd n77__vdd 62.5111
rk676 n73__vdd n78__vdd 62.4805
rk677 n76__vdd n79__vdd 77.78e-3
rk678 n79__vdd n1__vdd 85.67e-3
rk679 n1__vdd n80__vdd 100.1e-3
rk680 n80__vdd n81__vdd 15.8697
rk681 n76__vdd n82__vdd 62.5111
rk682 n80__vdd n83__vdd 100.9e-3
rk683 n83__vdd n84__vdd 15.8697
rk684 n80__vdd n85__vdd 15.8697
rk685 n83__vdd n86__vdd 276e-3
rk686 n86__vdd n87__vdd 62.5449
rk687 n83__vdd n88__vdd 15.8697
rk688 n86__vdd n89__vdd 30.6e-3
rk689 n89__vdd n90__vdd 277e-3
rk690 n90__vdd n91__vdd 31.2233
rk691 n86__vdd n92__vdd 62.5449
rk692 n90__vdd n93__vdd 31.2526
rk693 n16__vdd n17__vdd 5.3571
rk694 n16__vdd n25__vdd 3.75
rk695 n41__vdd n42__vdd 31
rk696 n55__vdd n56__vdd 31
rk697 n16__vdd n60__vdd 3.75
rk698 n16__vdd n79__vdd 3.75
rk699 n16__vdd n89__vdd 3.75
rk700 n47__vss n48__vss 37.7376
rk701 n48__vss n49__vss 50.46e-3
rk702 n49__vss n50__vss 64.12e-3
rk703 n50__vss n51__vss 37.03e-3
rk704 n51__vss n52__vss 27.09e-3
rk705 n52__vss n53__vss 74.05e-3
rk706 n53__vss n54__vss 26.87e-3
rk707 n54__vss n55__vss 31.84e-3
rk708 n55__vss n56__vss 50.46e-3
rk709 n56__vss n57__vss 50.46e-3
rk710 n57__vss n58__vss 101.4e-3
rk711 n58__vss n59__vss 101.4e-3
rk712 n59__vss n60__vss 39.51e-3
rk713 n60__vss n61__vss 25.85e-3
rk714 n61__vss n62__vss 40.53e-3
rk715 n62__vss n63__vss 78e-3
rk716 n63__vss n64__vss 23.37e-3
rk717 n64__vss n65__vss 24.39e-3
rk718 n65__vss n66__vss 39.29e-3
rk719 n66__vss n67__vss 113.3e-3
rk720 n67__vss n68__vss 12.68e-3
rk721 n68__vss n69__vss 165.9e-3
rk722 n69__vss n70__vss 69.31e-3
rk723 n70__vss n71__vss 55.65e-3
rk724 n71__vss vss 30.82e-3
rk725 vss n72__vss 85.63e-3
rk726 n72__vss n73__vss 61.82e-3
rk727 n73__vss n74__vss 54.19e-3
rk728 n74__vss n75__vss 46.74e-3
rk729 n75__vss n76__vss 16.94e-3
rk730 n76__vss n77__vss 65.36e-3
rk731 n77__vss n78__vss 35.56e-3
rk732 n78__vss n79__vss 82.74e-3
rk733 n79__vss n80__vss 55.65e-3
rk734 n80__vss n81__vss 186e-3
rk735 n81__vss n82__vss 101.4e-3
rk736 n82__vss n83__vss 16.94e-3
rk737 n83__vss n84__vss 46.74e-3
rk738 n84__vss n85__vss 54.19e-3
rk739 n85__vss n86__vss 61.82e-3
rk740 n86__vss n87__vss 125.4e-3
rk741 n48__vss n88__vss 37.6853
rk742 n49__vss n89__vss 37.6968
rk743 n50__vss n90__vss 37.6853
rk744 n51__vss n91__vss 37.6926
rk745 n52__vss n92__vss 37.6853
rk746 n53__vss n93__vss 37.691
rk747 n54__vss n94__vss 37.6853
rk748 n55__vss n95__vss 37.691
rk749 n56__vss n96__vss 75.2174
rk750 n57__vss n97__vss 37.6968
rk751 n58__vss n98__vss 37.6968
rk752 n59__vss n99__vss 37.6853
rk753 n61__vss n101__vss 219.9e-3
rk754 n62__vss n102__vss 37.6853
rk755 n64__vss n103__vss 37.6853
rk756 n65__vss n104__vss 37.6983
rk757 n66__vss n105__vss 75.222
rk758 n67__vss n106__vss 75.2251
rk759 n68__vss n107__vss 37.6983
rk760 n69__vss n109__vss 222e-3
rk761 n109__vss n110__vss 31.4165
rk762 n71__vss n111__vss 37.6853
rk763 n72__vss n112__vss 37.7565
rk764 n72__vss n113__vss 37.7592
rk765 n73__vss n114__vss 37.6853
rk766 n74__vss n115__vss 37.6853
rk767 n75__vss n116__vss 37.6853
rk768 n76__vss n117__vss 37.6853
rk769 n77__vss n118__vss 75.2174
rk770 n78__vss n119__vss 37.6853
rk771 n79__vss n120__vss 75.2174
rk772 n81__vss n121__vss 37.6853
rk773 n82__vss n122__vss 37.6853
rk774 n83__vss n123__vss 37.6853
rk775 n84__vss n124__vss 75.222
rk776 n85__vss n125__vss 37.6853
rk777 n86__vss n126__vss 75.2932
rk778 n86__vss n127__vss 75.2935
rk779 n87__vss n128__vss 75.2154
rk780 n87__vss n129__vss 75.4156
rk781 n101__vss n130__vss 31.4157
rk782 n3__vss n51__vss 4.4286
rk783 n3__vss n60__vss 3.1
rk784 n3__vss n70__vss 3.1
rk785 n3__vss n80__vss 3.1
rk786 n3__vss n87__vss 3.1
rk787 n100__vss n101__vss 75
rk788 n108__vss n109__vss 75
rk789 n94__vdd n95__vdd 15.8453
rk790 n95__vdd n96__vdd 107.7e-3
rk791 n96__vdd n98__vdd 36.81e-3
rk792 n98__vdd n99__vdd 26.87e-3
rk793 n99__vdd n100__vdd 100.9e-3
rk794 n100__vdd n101__vdd 114.6e-3
rk795 n101__vdd n102__vdd 63.68e-3
rk796 n102__vdd n103__vdd 197e-3
rk797 n103__vdd n104__vdd 66.6e-3
rk798 n104__vdd n105__vdd 100.9e-3
rk799 n105__vdd n106__vdd 276e-3
rk800 n106__vdd n107__vdd 149.8e-3
rk801 n107__vdd vdd 86.91e-3
rk802 vdd n108__vdd 87.71e-3
rk803 n108__vdd n109__vdd 114.6e-3
rk804 n109__vdd n110__vdd 63.68e-3
rk805 n110__vdd n111__vdd 100.9e-3
rk806 n111__vdd n112__vdd 114.6e-3
rk807 n112__vdd n113__vdd 23.15e-3
rk808 n113__vdd n4__vdd 85.67e-3
rk809 n95__vdd n114__vdd 15.7861
rk810 n96__vdd n115__vdd 15.8697
rk811 n96__vdd n116__vdd 15.8697
rk812 n99__vdd n117__vdd 15.8697
rk813 n99__vdd n118__vdd 15.8697
rk814 n100__vdd n119__vdd 15.8697
rk815 n100__vdd n120__vdd 15.8697
rk816 n101__vdd n121__vdd 62.4805
rk817 n101__vdd n122__vdd 62.4805
rk818 n102__vdd n123__vdd 62.5111
rk819 n102__vdd n124__vdd 62.5111
rk820 n104__vdd n125__vdd 15.8697
rk821 n104__vdd n126__vdd 15.8697
rk822 n105__vdd n127__vdd 15.8697
rk823 n105__vdd n128__vdd 15.8697
rk824 n106__vdd n129__vdd 62.5449
rk825 n106__vdd n130__vdd 62.5449
rk826 n108__vdd n131__vdd 15.8697
rk827 n108__vdd n132__vdd 15.8697
rk828 n109__vdd n133__vdd 15.8697
rk829 n109__vdd n134__vdd 15.8697
rk830 n110__vdd n135__vdd 15.8697
rk831 n110__vdd n136__vdd 15.8697
rk832 n111__vdd n137__vdd 15.8697
rk833 n111__vdd n138__vdd 15.8697
rk834 n112__vdd n139__vdd 62.4805
rk835 n112__vdd n140__vdd 62.4805
rk836 n4__vdd n141__vdd 62.4142
rk837 n4__vdd n142__vdd 219.3e-3
rk838 n142__vdd n143__vdd 15.8697
rk839 n4__vdd n144__vdd 62.4142
rk840 n142__vdd n145__vdd 100.9e-3
rk841 n145__vdd n146__vdd 15.8697
rk842 n142__vdd n147__vdd 15.8697
rk843 n145__vdd n148__vdd 188.3e-3
rk844 n148__vdd n149__vdd 87.71e-3
rk845 n149__vdd n150__vdd 62.5449
rk846 n145__vdd n151__vdd 15.8697
rk848 n149__vdd n153__vdd 62.5449
rk849 n97__vdd n98__vdd 5.3571
rk850 n97__vdd n103__vdd 3.75
rk851 n97__vdd n107__vdd 3.75
rk852 n97__vdd n113__vdd 3.75
rk853 n97__vdd n148__vdd 3.75
rk854 n131__vss n132__vss 37.7536
rk855 n132__vss n133__vss 107.7e-3
rk856 n133__vss n134__vss 36.81e-3
rk857 n134__vss n135__vss 26.87e-3
rk858 n135__vss n136__vss 100.9e-3
rk859 n136__vss n137__vss 82.3e-3
rk860 n137__vss n138__vss 293.8e-3
rk861 n138__vss n139__vss 66.6e-3
rk862 n139__vss n140__vss 77.78e-3
rk863 n140__vss n141__vss 23.15e-3
rk864 n141__vss n142__vss 63.68e-3
rk865 n142__vss n143__vss 114.6e-3
rk866 n143__vss n144__vss 246.6e-3
rk867 n144__vss vss 86.91e-3
rk868 vss n145__vss 87.71e-3
rk869 n145__vss n146__vss 114.6e-3
rk870 n146__vss n147__vss 63.68e-3
rk871 n147__vss n148__vss 100.9e-3
rk872 n148__vss n149__vss 82.3e-3
rk873 n149__vss n150__vss 55.43e-3
rk874 n150__vss n151__vss 305e-3
rk875 n151__vss n152__vss 100.9e-3
rk876 n152__vss n153__vss 63.68e-3
rk877 n153__vss n154__vss 123.7e-3
rk878 n132__vss n155__vss 37.6944
rk879 n133__vss n156__vss 37.778
rk880 n133__vss n157__vss 37.778
rk881 n135__vss n158__vss 37.778
rk882 n135__vss n159__vss 37.778
rk883 n136__vss n160__vss 37.778
rk884 n136__vss n161__vss 37.778
rk885 n137__vss n162__vss 75.3101
rk886 n137__vss n163__vss 75.3101
rk887 n139__vss n164__vss 37.778
rk888 n139__vss n165__vss 37.778
rk889 n141__vss n166__vss 37.778
rk890 n141__vss n167__vss 37.778
rk891 n142__vss n168__vss 75.3147
rk892 n142__vss n169__vss 75.3147
rk893 n143__vss n170__vss 75.3123
rk894 n143__vss n171__vss 75.3123
rk895 n145__vss n172__vss 37.778
rk896 n145__vss n173__vss 37.778
rk897 n146__vss n174__vss 37.778
rk898 n146__vss n175__vss 37.778
rk899 n147__vss n176__vss 37.778
rk900 n147__vss n177__vss 37.778
rk901 n148__vss n178__vss 37.778
rk902 n148__vss n179__vss 37.778
rk903 n149__vss n180__vss 75.3101
rk904 n149__vss n181__vss 75.3101
rk905 n151__vss n182__vss 37.778
rk906 n151__vss n183__vss 37.778
rk907 n152__vss n184__vss 37.778
rk908 n152__vss n185__vss 37.778
rk909 n153__vss n186__vss 75.3147
rk910 n153__vss n187__vss 75.3147
rk911 n154__vss n188__vss 75.2154
rk912 n154__vss n189__vss 75.2154
rk913 n3__vss n134__vss 4.4286
rk914 n3__vss n138__vss 3.1
rk915 n3__vss n144__vss 3.1
rk916 n3__vss n150__vss 3.1
rk917 n3__vss n154__vss 3.1
rk918 n154__vdd n155__vdd 15.8453
rk919 n155__vdd n156__vdd 107.7e-3
rk920 n156__vdd n158__vdd 36.81e-3
rk921 n158__vdd n159__vdd 26.87e-3
rk922 n159__vdd n160__vdd 100.9e-3
rk923 n160__vdd n161__vdd 114.6e-3
rk924 n161__vdd n162__vdd 63.68e-3
rk925 n162__vdd n163__vdd 197e-3
rk926 n163__vdd n164__vdd 66.6e-3
rk927 n164__vdd n165__vdd 100.9e-3
rk928 n165__vdd n166__vdd 276e-3
rk929 n166__vdd n167__vdd 149.8e-3
rk930 n167__vdd vdd 86.91e-3
rk931 vdd n168__vdd 87.71e-3
rk932 n168__vdd n169__vdd 114.6e-3
rk933 n169__vdd n170__vdd 63.68e-3
rk934 n170__vdd n171__vdd 100.9e-3
rk935 n171__vdd n172__vdd 114.6e-3
rk936 n172__vdd n173__vdd 23.15e-3
rk937 n173__vdd n5__vdd 85.67e-3
rk938 n155__vdd n174__vdd 15.7861
rk939 n156__vdd n175__vdd 15.8697
rk940 n156__vdd n176__vdd 15.8697
rk941 n159__vdd n177__vdd 15.8697
rk942 n159__vdd n178__vdd 15.8697
rk943 n160__vdd n179__vdd 15.8697
rk944 n160__vdd n180__vdd 15.8697
rk945 n161__vdd n181__vdd 62.4805
rk946 n161__vdd n182__vdd 62.4805
rk947 n162__vdd n183__vdd 62.5111
rk948 n162__vdd n184__vdd 62.5111
rk949 n164__vdd n185__vdd 15.8697
rk950 n164__vdd n186__vdd 15.8697
rk951 n165__vdd n187__vdd 15.8697
rk952 n165__vdd n188__vdd 15.8697
rk953 n166__vdd n189__vdd 62.5449
rk954 n166__vdd n190__vdd 62.5449
rk955 n168__vdd n191__vdd 15.8697
rk956 n168__vdd n192__vdd 15.8697
rk957 n169__vdd n193__vdd 15.8697
rk958 n169__vdd n194__vdd 15.8697
rk959 n170__vdd n195__vdd 15.8697
rk960 n170__vdd n196__vdd 15.8697
rk961 n171__vdd n197__vdd 15.8697
rk962 n171__vdd n198__vdd 15.8697
rk963 n172__vdd n199__vdd 62.4805
rk964 n172__vdd n200__vdd 62.4805
rk965 n5__vdd n201__vdd 62.4142
rk966 n5__vdd n202__vdd 219.3e-3
rk967 n202__vdd n203__vdd 15.8697
rk968 n5__vdd n204__vdd 62.4142
rk969 n202__vdd n205__vdd 100.9e-3
rk970 n205__vdd n206__vdd 15.8697
rk971 n202__vdd n207__vdd 15.8697
rk972 n205__vdd n208__vdd 188.3e-3
rk973 n208__vdd n209__vdd 87.71e-3
rk974 n209__vdd n210__vdd 62.5449
rk975 n205__vdd n211__vdd 15.8697
rk977 n209__vdd n213__vdd 62.5449
rk978 n157__vdd n158__vdd 5.3571
rk979 n157__vdd n163__vdd 3.75
rk980 n157__vdd n167__vdd 3.75
rk981 n157__vdd n173__vdd 3.75
rk982 n157__vdd n208__vdd 3.75
rk983 n190__vss n191__vss 37.8034
rk984 n191__vss n192__vss 37.03e-3
rk985 n192__vss n193__vss 27.09e-3
rk986 n193__vss n194__vss 101.4e-3
rk987 n194__vss n195__vss 82.74e-3
rk988 n195__vss n196__vss 294e-3
rk989 n196__vss n197__vss 66.82e-3
rk990 n197__vss n198__vss 78e-3
rk991 n198__vss n199__vss 23.37e-3
rk992 n199__vss n200__vss 64.12e-3
rk993 n200__vss n201__vss 115e-3
rk994 n201__vss n202__vss 246.8e-3
rk995 n202__vss vss 86.91e-3
rk996 vss n203__vss 87.93e-3
rk997 n203__vss n204__vss 115e-3
rk998 n204__vss n205__vss 64.12e-3
rk999 n205__vss n206__vss 101.4e-3
rk1000 n206__vss n207__vss 82.74e-3
rk1001 n207__vss n208__vss 55.65e-3
rk1002 n208__vss n209__vss 305.2e-3
rk1003 n209__vss n210__vss 101.4e-3
rk1004 n210__vss n211__vss 64.12e-3
rk1005 n211__vss n212__vss 123.9e-3
rk1006 n191__vss n213__vss 37.6853
rk1007 n193__vss n214__vss 37.6853
rk1008 n194__vss n215__vss 37.6853
rk1009 n195__vss n216__vss 75.2174
rk1010 n197__vss n217__vss 37.6853
rk1011 n199__vss n218__vss 37.6853
rk1012 n200__vss n219__vss 75.222
rk1013 n201__vss n220__vss 75.2196
rk1014 n203__vss n221__vss 37.6853
rk1015 n204__vss n222__vss 37.6853
rk1016 n205__vss n223__vss 37.6853
rk1017 n206__vss n224__vss 37.6853
rk1018 n207__vss n225__vss 75.2174
rk1019 n209__vss n226__vss 37.6853
rk1020 n210__vss n227__vss 37.6853
rk1021 n211__vss n228__vss 75.222
rk1022 n212__vss n229__vss 75.2154
rk1023 n3__vss n192__vss 4.4286
rk1024 n3__vss n196__vss 3.1
rk1025 n3__vss n202__vss 3.1
rk1026 n3__vss n208__vss 3.1
rk1027 n3__vss n212__vss 3.1
rl1 n1__clk n2__clk 202.615
rl2 n2__clk n3__clk 33.3841
rl3 n1__rst n2__rst 152.615
rl4 n2__rst n3__rst 83.3841
rl5 net9 n2__net9 126.36
rl6 net10 n2__net10 87.898
rl7 n3__net10 n4__net10 87.898
rl8 n3__net9 n4__net9 126.36
rl9 n5__net9 n6__net9 126.36
rl10 n5__net10 n6__net10 87.898
rl11 n7__net10 n8__net10 87.898
rl12 n7__net9 n8__net9 126.36
rl13 i0__net3 n2__i0__net3 126.36
rl14 n4__clk n5__clk 87.898
rl15 i0__net7 n2__i0__net7 87.898
rl16 i0__net1 n2__i0__net1 126.36
rl17 i1__net2 n2__i1__net2 11.2742
rl18 i1__net2 n3__i1__net2 9.7184
rl19 i2__net2 n2__i2__net2 9.7184
rl20 i2__net2 n3__i2__net2 11.2742
rl21 i3__net2 n2__i3__net2 11.2742
rl22 i3__net2 n3__i3__net2 9.7184
rl23 i8__net2 n2__i8__net2 9.7184
rl24 i8__net2 n3__i8__net2 11.2742
rl25 i0__i2__net2 n2__i0__i2__net2 11.2742
rl26 i0__i2__net2 n3__i0__i2__net2 9.7184
rl27 i0__i3__net2 n2__i0__i3__net2 9.7184
rl28 i0__i3__net2 n3__i0__i3__net2 11.2742
rl29 net3 n2__net3 98.1035
rl30 n3__net3 n4__net3 98.1035
rl31 n5__net3 n6__net3 98.1035
rl32 n7__net3 n8__net3 98.1035
rl33 n4__rst n5__rst 98.1035
rl34 n6__rst n7__rst 98.1035
rl35 i1__net1 n2__i1__net1 56.5719
rl36 n2__i1__net1 n3__i1__net1 23.6889
rl37 n3__i1__net1 n4__i1__net1 50.6296
rl38 n2__i1__net1 n5__i1__net1 56.5719
rl39 n3__i1__net1 n6__i1__net1 55.6157
rl40 n3__i1__net1 n7__i1__net1 55.6157
rl41 i2__net1 n2__i2__net1 56.5719
rl42 n2__i2__net1 n3__i2__net1 23.6889
rl43 n3__i2__net1 n4__i2__net1 50.6296
rl44 n2__i2__net1 n5__i2__net1 56.5719
rl45 n3__i2__net1 n6__i2__net1 55.6157
rl46 n3__i2__net1 n7__i2__net1 55.6157
rl47 i3__net1 n2__i3__net1 56.5719
rl48 n2__i3__net1 n3__i3__net1 23.6889
rl49 n3__i3__net1 n4__i3__net1 50.6296
rl50 n2__i3__net1 n5__i3__net1 56.5719
rl51 n3__i3__net1 n6__i3__net1 55.6157
rl52 n3__i3__net1 n7__i3__net1 55.6157
rl53 i8__net1 n2__i8__net1 56.5719
rl54 n2__i8__net1 n3__i8__net1 23.6889
rl55 n3__i8__net1 n4__i8__net1 50.6296
rl56 n2__i8__net1 n5__i8__net1 56.5719
rl57 n3__i8__net1 n6__i8__net1 55.6157
rl58 n3__i8__net1 n7__i8__net1 55.6157
rl59 i0__i2__net1 n2__i0__i2__net1 56.5719
rl60 n2__i0__i2__net1 n3__i0__i2__net1 23.6889
rl61 n3__i0__i2__net1 n4__i0__i2__net1 50.6296
rl62 n2__i0__i2__net1 n5__i0__i2__net1 56.5719
rl63 n3__i0__i2__net1 n6__i0__i2__net1 55.6157
rl64 n3__i0__i2__net1 n7__i0__i2__net1 55.6157
rl65 i0__i3__net1 n2__i0__i3__net1 56.5719
rl66 n2__i0__i3__net1 n3__i0__i3__net1 23.6889
rl67 n3__i0__i3__net1 n4__i0__i3__net1 50.6296
rl68 n2__i0__i3__net1 n5__i0__i3__net1 56.5719
rl69 n3__i0__i3__net1 n6__i0__i3__net1 55.6157
rl70 n3__i0__i3__net1 n7__i0__i3__net1 55.6157
rl71 n9__net10 n10__net10 126.36
rl72 n9__net9 n10__net9 87.898
rl73 n11__net9 n12__net9 87.898
rl74 n11__net10 n12__net10 126.36
rl75 n13__net10 n14__net10 126.36
rl76 n13__net9 n14__net9 87.898
rl77 n15__net9 n16__net9 87.898
rl78 n15__net10 n16__net10 126.36
rl79 n6__clk n7__clk 126.36
rl80 n3__i0__net3 n4__i0__net3 87.898
rl81 n3__i0__net1 n4__i0__net1 87.898
rl82 n3__i0__net7 n4__i0__net7 126.36
rl83 i1__net4 n2__i1__net4 11.2742
rl84 i1__net4 n3__i1__net4 9.7184
rl85 i2__net4 n2__i2__net4 9.7184
rl86 i2__net4 n3__i2__net4 11.2742
rl87 i3__net4 n2__i3__net4 11.2742
rl88 i3__net4 n3__i3__net4 9.7184
rl89 i8__net4 n2__i8__net4 9.7184
rl90 i8__net4 n3__i8__net4 11.2742
rl91 net4 n2__net4 74.5009
rl92 n3__net4 n4__net4 74.5009
rl93 n5__net4 n6__net4 74.5009
rl94 n7__net4 n8__net4 74.5009
rl95 i0__i2__net4 n2__i0__i2__net4 11.2742
rl96 i0__i2__net4 n3__i0__i2__net4 9.7184
rl97 i0__i3__net4 n2__i0__i3__net4 9.7184
rl98 i0__i3__net4 n3__i0__i3__net4 11.2742
rl99 i0__net6 n2__i0__net6 74.5009
rl100 n3__i0__net6 n4__i0__net6 74.5009
rl101 i1__net5 n2__i1__net5 56.5719
rl102 n2__i1__net5 n3__i1__net5 23.6889
rl103 n3__i1__net5 n4__i1__net5 50.6296
rl104 n2__i1__net5 n5__i1__net5 56.5719
rl105 n3__i1__net5 n6__i1__net5 55.6157
rl106 n3__i1__net5 n7__i1__net5 55.6157
rl107 i2__net5 n2__i2__net5 56.5719
rl108 n2__i2__net5 n3__i2__net5 23.6889
rl109 n3__i2__net5 n4__i2__net5 50.6296
rl110 n2__i2__net5 n5__i2__net5 56.5719
rl111 n3__i2__net5 n6__i2__net5 55.6157
rl112 n3__i2__net5 n7__i2__net5 55.6157
rl113 i3__net5 n2__i3__net5 56.5719
rl114 n2__i3__net5 n3__i3__net5 23.6889
rl115 n3__i3__net5 n4__i3__net5 50.6296
rl116 n2__i3__net5 n5__i3__net5 56.5719
rl117 n3__i3__net5 n6__i3__net5 55.6157
rl118 n3__i3__net5 n7__i3__net5 55.6157
rl119 i8__net5 n2__i8__net5 56.5719
rl120 n2__i8__net5 n3__i8__net5 23.6889
rl121 n3__i8__net5 n4__i8__net5 50.6296
rl122 n2__i8__net5 n5__i8__net5 56.5719
rl123 n3__i8__net5 n6__i8__net5 55.6157
rl124 n3__i8__net5 n7__i8__net5 55.6157
rl125 n4__i1__net4 n5__i1__net4 49.0903
rl126 n5__i1__net4 n6__i1__net4 49.0903
rl127 n4__i2__net4 n5__i2__net4 49.0903
rl128 n5__i2__net4 n6__i2__net4 49.0903
rl129 n4__i3__net4 n5__i3__net4 49.0903
rl130 n5__i3__net4 n6__i3__net4 49.0903
rl131 n4__i8__net4 n5__i8__net4 49.0903
rl132 n5__i8__net4 n6__i8__net4 49.0903
rl133 i0__i2__net5 n2__i0__i2__net5 56.5719
rl134 n2__i0__i2__net5 n3__i0__i2__net5 23.6889
rl135 n3__i0__i2__net5 n4__i0__i2__net5 50.6296
rl136 n2__i0__i2__net5 n5__i0__i2__net5 56.5719
rl137 n3__i0__i2__net5 n6__i0__i2__net5 55.6157
rl138 n3__i0__i2__net5 n7__i0__i2__net5 55.6157
rl139 i0__i3__net5 n2__i0__i3__net5 56.5719
rl140 n2__i0__i3__net5 n3__i0__i3__net5 23.6889
rl141 n3__i0__i3__net5 n4__i0__i3__net5 50.6296
rl142 n2__i0__i3__net5 n5__i0__i3__net5 56.5719
rl143 n3__i0__i3__net5 n6__i0__i3__net5 55.6157
rl144 n3__i0__i3__net5 n7__i0__i3__net5 55.6157
rl145 n1__x_out_b_3 n2__x_out_b_3 56.5719
rl146 n2__x_out_b_3 n3__x_out_b_3 50.013
rl147 n2__x_out_b_3 n4__x_out_b_3 56.5719
rl148 n1__x_out_b_2 n2__x_out_b_2 56.5719
rl149 n2__x_out_b_2 n3__x_out_b_2 50.013
rl150 n2__x_out_b_2 n4__x_out_b_2 56.5719
rl151 n1__x_out_b_1 n2__x_out_b_1 56.5719
rl152 n2__x_out_b_1 n3__x_out_b_1 50.013
rl153 n2__x_out_b_1 n4__x_out_b_1 56.5719
rl154 n1__x_out_b_0 n2__x_out_b_0 56.5719
rl155 n2__x_out_b_0 n3__x_out_b_0 50.013
rl156 n2__x_out_b_0 n4__x_out_b_0 56.5719
rl157 n4__i0__i2__net4 n5__i0__i2__net4 49.0903
rl158 n5__i0__i2__net4 n6__i0__i2__net4 49.0903
rl159 n4__i0__i3__net4 n5__i0__i3__net4 49.0903
rl160 n5__i0__i3__net4 n6__i0__i3__net4 49.0903
rl161 n14__i0__net1 n15__i0__net1 56.5719
rl162 n15__i0__net1 n16__i0__net1 50.013
rl163 n15__i0__net1 n17__i0__net1 56.5719
rl164 n6__i0__net8 n7__i0__net8 56.5719
rl165 n7__i0__net8 n8__i0__net8 50.013
rl166 n7__i0__net8 n9__i0__net8 56.5719
rl167 n33__net9 n34__net9 126.36
rl168 n41__net10 n42__net10 87.898
rl169 n43__net10 n44__net10 87.898
rl170 n35__net9 n36__net9 126.36
rl171 n37__net9 n38__net9 126.36
rl172 n45__net10 n46__net10 87.898
rl173 n47__net10 n48__net10 87.898
rl174 n39__net9 n40__net9 126.36
rl175 i0__net10 n2__i0__net10 56.5719
rl176 n2__i0__net10 n3__i0__net10 48.1183
rl177 n2__i0__net10 n4__i0__net10 56.5719
rl178 n10__i0__net8 n11__i0__net8 69.2328
rl179 i0__net11 n2__i0__net11 101.925
rl180 n2__i0__net11 n3__i0__net11 201.489
rl181 n12__i0__net8 n13__i0__net8 73.079
rl182 i0__net9 n2__i0__net9 56.5719
rl183 n2__i0__net9 n3__i0__net9 48.1183
rl184 n2__i0__net9 n4__i0__net9 56.5719
rl185 i7__net2 n2__i7__net2 11.2742
rl186 i7__net2 n3__i7__net2 9.7184
rl187 i6__net2 n2__i6__net2 9.7184
rl188 i6__net2 n3__i6__net2 11.2742
rl189 i4__net2 n2__i4__net2 11.2742
rl190 i4__net2 n3__i4__net2 9.7184
rl191 i5__net2 n2__i5__net2 9.7184
rl192 i5__net2 n3__i5__net2 11.2742
rl193 n5__i0__net9 n6__i0__net9 64.1533
rl194 n6__i0__net9 n7__i0__net9 33.3841
rl195 n29__net3 n30__net3 98.1035
rl196 n31__net3 n32__net3 98.1035
rl197 n33__net3 n34__net3 98.1035
rl198 n35__net3 n36__net3 98.1035
rl199 n5__i0__net10 n6__i0__net10 33.3841
rl200 n6__i0__net10 n7__i0__net10 64.1533
rl201 n4__i0__net11 n5__i0__net11 73.079
rl202 i7__net1 n2__i7__net1 56.5719
rl203 n2__i7__net1 n3__i7__net1 23.6889
rl204 n3__i7__net1 n4__i7__net1 50.6296
rl205 n2__i7__net1 n5__i7__net1 56.5719
rl206 n3__i7__net1 n6__i7__net1 55.6157
rl207 n3__i7__net1 n7__i7__net1 55.6157
rl208 i6__net1 n2__i6__net1 56.5719
rl209 n2__i6__net1 n3__i6__net1 23.6889
rl210 n3__i6__net1 n4__i6__net1 50.6296
rl211 n2__i6__net1 n5__i6__net1 56.5719
rl212 n3__i6__net1 n6__i6__net1 55.6157
rl213 n3__i6__net1 n7__i6__net1 55.6157
rl214 i4__net1 n2__i4__net1 56.5719
rl215 n2__i4__net1 n3__i4__net1 23.6889
rl216 n3__i4__net1 n4__i4__net1 50.6296
rl217 n2__i4__net1 n5__i4__net1 56.5719
rl218 n3__i4__net1 n6__i4__net1 55.6157
rl219 n3__i4__net1 n7__i4__net1 55.6157
rl220 i5__net1 n2__i5__net1 56.5719
rl221 n2__i5__net1 n3__i5__net1 23.6889
rl222 n3__i5__net1 n4__i5__net1 50.6296
rl223 n2__i5__net1 n5__i5__net1 56.5719
rl224 n3__i5__net1 n6__i5__net1 55.6157
rl225 n3__i5__net1 n7__i5__net1 55.6157
rl226 n14__i0__net8 n15__i0__net8 201.489
rl227 n15__i0__net8 n16__i0__net8 69.2328
rl228 n6__i0__net11 n7__i0__net11 101.925
rl229 n23__rst n24__rst 56.5719
rl230 n24__rst n25__rst 23.6889
rl231 n25__rst n26__rst 10.1559
rl232 n26__rst n27__rst 8.8401
rl233 n27__rst n28__rst 26.2002
rl234 n28__rst n29__rst 9.498
rl235 n29__rst n30__rst 9.498
rl236 n30__rst n31__rst 23.6922
rl237 n31__rst n32__rst 56.5719
rl238 n24__rst n33__rst 56.5719
rl239 n25__rst n34__rst 55.6157
rl240 n25__rst n35__rst 55.6157
rl241 n27__rst n36__rst 55.6157
rl242 n27__rst n37__rst 55.6157
rl243 n28__rst n38__rst 55.6157
rl244 n28__rst n39__rst 55.6157
rl245 n30__rst n40__rst 55.6157
rl246 n30__rst n41__rst 55.6157
rl247 n31__rst n42__rst 56.5719
rl248 n57__net10 n58__net10 126.36
rl249 n49__net9 n50__net9 87.898
rl250 n51__net9 n52__net9 87.898
rl251 n59__net10 n60__net10 126.36
rl252 n61__net10 n62__net10 126.36
rl253 n53__net9 n54__net9 87.898
rl254 n55__net9 n56__net9 87.898
rl255 n63__net10 n64__net10 126.36
rl256 net7 n2__net7 56.5719
rl257 n2__net7 n3__net7 48.1183
rl258 n2__net7 n4__net7 56.5719
rl259 i7__net4 n2__i7__net4 11.2742
rl260 i7__net4 n3__i7__net4 9.7184
rl261 i6__net4 n2__i6__net4 9.7184
rl262 i6__net4 n3__i6__net4 11.2742
rl263 i4__net4 n2__i4__net4 11.2742
rl264 i4__net4 n3__i4__net4 9.7184
rl265 i5__net4 n2__i5__net4 9.7184
rl266 i5__net4 n3__i5__net4 11.2742
rl267 n21__net4 n22__net4 74.5009
rl268 n23__net4 n24__net4 74.5009
rl269 n25__net4 n26__net4 74.5009
rl270 n27__net4 n28__net4 74.5009
rl271 net11 n2__net11 56.5719
rl272 n2__net11 n3__net11 48.1183
rl273 n2__net11 n4__net11 56.5719
rl274 n29__net4 n30__net4 56.5719
rl275 n30__net4 n31__net4 23.6889
rl276 n31__net4 n32__net4 9.498
rl277 n32__net4 n33__net4 9.498
rl278 n33__net4 n34__net4 26.2002
rl279 n34__net4 n35__net4 9.498
rl280 n35__net4 n36__net4 9.498
rl281 n36__net4 n37__net4 23.6922
rl282 n37__net4 n38__net4 56.5719
rl283 n30__net4 n39__net4 56.5719
rl284 n31__net4 n40__net4 55.6157
rl285 n31__net4 n41__net4 55.6157
rl286 n33__net4 n42__net4 55.6157
rl287 n33__net4 n43__net4 55.6157
rl288 n34__net4 n44__net4 55.6157
rl289 n34__net4 n45__net4 55.6157
rl290 n36__net4 n46__net4 55.6157
rl291 n36__net4 n47__net4 55.6157
rl292 n37__net4 n48__net4 56.5719
rl293 i7__net5 n2__i7__net5 56.5719
rl294 n2__i7__net5 n3__i7__net5 23.6889
rl295 n3__i7__net5 n4__i7__net5 50.6296
rl296 n2__i7__net5 n5__i7__net5 56.5719
rl297 n3__i7__net5 n6__i7__net5 55.6157
rl298 n3__i7__net5 n7__i7__net5 55.6157
rl299 i6__net5 n2__i6__net5 56.5719
rl300 n2__i6__net5 n3__i6__net5 23.6889
rl301 n3__i6__net5 n4__i6__net5 50.6296
rl302 n2__i6__net5 n5__i6__net5 56.5719
rl303 n3__i6__net5 n6__i6__net5 55.6157
rl304 n3__i6__net5 n7__i6__net5 55.6157
rl305 i4__net5 n2__i4__net5 56.5719
rl306 n2__i4__net5 n3__i4__net5 23.6889
rl307 n3__i4__net5 n4__i4__net5 50.6296
rl308 n2__i4__net5 n5__i4__net5 56.5719
rl309 n3__i4__net5 n6__i4__net5 55.6157
rl310 n3__i4__net5 n7__i4__net5 55.6157
rl311 i5__net5 n2__i5__net5 56.5719
rl312 n2__i5__net5 n3__i5__net5 23.6889
rl313 n3__i5__net5 n4__i5__net5 50.6296
rl314 n2__i5__net5 n5__i5__net5 56.5719
rl315 n3__i5__net5 n6__i5__net5 55.6157
rl316 n3__i5__net5 n7__i5__net5 55.6157
rl317 n4__i7__net4 n5__i7__net4 49.0903
rl318 n5__i7__net4 n6__i7__net4 49.0903
rl319 n4__i6__net4 n5__i6__net4 49.0903
rl320 n5__i6__net4 n6__i6__net4 49.0903
rl321 n4__i4__net4 n5__i4__net4 49.0903
rl322 n5__i4__net4 n6__i4__net4 49.0903
rl323 n4__i5__net4 n5__i5__net4 49.0903
rl324 n5__i5__net4 n6__i5__net4 49.0903
rl325 n5__net7 n6__net7 56.5719
rl326 n6__net7 n7__net7 23.6889
rl327 n7__net7 n8__net7 9.498
rl328 n8__net7 n9__net7 9.498
rl329 n9__net7 n10__net7 26.2002
rl330 n10__net7 n11__net7 9.498
rl331 n11__net7 n12__net7 9.498
rl332 n12__net7 n13__net7 23.6922
rl333 n13__net7 n14__net7 56.5719
rl334 n6__net7 n15__net7 56.5719
rl335 n7__net7 n16__net7 55.6157
rl336 n7__net7 n17__net7 55.6157
rl337 n9__net7 n18__net7 55.6157
rl338 n9__net7 n19__net7 55.6157
rl339 n10__net7 n20__net7 55.6157
rl340 n10__net7 n21__net7 55.6157
rl341 n12__net7 n22__net7 55.6157
rl342 n12__net7 n23__net7 55.6157
rl343 n13__net7 n24__net7 56.5719
rl344 n5__net11 n6__net11 56.5719
rl345 n6__net11 n7__net11 23.6889
rl346 n7__net11 n8__net11 9.498
rl347 n8__net11 n9__net11 9.498
rl348 n9__net11 n10__net11 26.2002
rl349 n10__net11 n11__net11 9.498
rl350 n11__net11 n12__net11 9.498
rl351 n12__net11 n13__net11 23.6922
rl352 n13__net11 n14__net11 56.5719
rl353 n6__net11 n15__net11 56.5719
rl354 n7__net11 n16__net11 55.6157
rl355 n7__net11 n17__net11 55.6157
rl356 n9__net11 n18__net11 55.6157
rl357 n9__net11 n19__net11 55.6157
rl358 n10__net11 n20__net11 55.6157
rl359 n10__net11 n21__net11 55.6157
rl360 n12__net11 n22__net11 55.6157
rl361 n12__net11 n23__net11 55.6157
rl362 n13__net11 n24__net11 56.5719
rl363 n1__y_out_b_3 n2__y_out_b_3 56.5719
rl364 n2__y_out_b_3 n3__y_out_b_3 50.013
rl365 n2__y_out_b_3 n4__y_out_b_3 56.5719
rl366 n1__y_out_b_2 n2__y_out_b_2 56.5719
rl367 n2__y_out_b_2 n3__y_out_b_2 50.013
rl368 n2__y_out_b_2 n4__y_out_b_2 56.5719
rl369 n1__y_out_b_1 n2__y_out_b_1 56.5719
rl370 n2__y_out_b_1 n3__y_out_b_1 50.013
rl371 n2__y_out_b_1 n4__y_out_b_1 56.5719
rl372 n1__y_out_b_0 n2__y_out_b_0 56.5719
rl373 n2__y_out_b_0 n3__y_out_b_0 50.013
rl374 n2__y_out_b_0 n4__y_out_b_0 56.5719
mpm2_5__rcx n30__vdd n22__net7 n75__net9 n16__vdd g45p1svt L=45e-9 W=480e-9 AD=76.8e-15 AS=76.8e-15 PD=1.28e-6 PS=1.28e-6 NRD=1.16667 NRS=1.16667 M=1
mpm2_4__rcx n78__net9 n20__net7 n30__vdd n16__vdd g45p1svt L=45e-9 W=480e-9 AD=76.8e-15 AS=76.8e-15 PD=1.28e-6 PS=1.28e-6 NRD=1.16667 NRS=1.16667 M=1
mpm2_3__rcx n28__vdd n18__net7 n78__net9 n16__vdd g45p1svt L=45e-9 W=480e-9 AD=76.8e-15 AS=76.8e-15 PD=1.28e-6 PS=1.28e-6 NRD=1.16667 NRS=1.16667 M=1
mpm2_2__rcx n81__net9 n16__net7 n28__vdd n16__vdd g45p1svt L=45e-9 W=480e-9 AD=76.8e-15 AS=76.8e-15 PD=1.28e-6 PS=1.28e-6 NRD=1.16667 NRS=1.16667 M=1
mpm2_1__rcx n13__vdd n15__net7 n81__net9 n16__vdd g45p1svt L=45e-9 W=480e-9 AD=67.2e-15 AS=67.2e-15 PD=1.26e-6 PS=1.26e-6 NRD=1.16667 NRS=1.16667 M=1
mpm2 n75__net9 n14__net7 n32__vdd n16__vdd g45p1svt L=45e-9 W=480e-9 AD=76.8e-15 AS=76.8e-15 PD=1.26e-6 PS=1.26e-6 NRD=1.16667 NRS=1.16667 M=1
mpm8_5__rcx n51__vdd n40__rst n51__net4 n16__vdd g45p1svt L=45e-9 W=480e-9 AD=76.8e-15 AS=76.8e-15 PD=1.28e-6 PS=1.28e-6 NRD=1.16667 NRS=1.16667 M=1
mpm8_4__rcx n54__net4 n38__rst n51__vdd n16__vdd g45p1svt L=45e-9 W=480e-9 AD=76.8e-15 AS=76.8e-15 PD=1.28e-6 PS=1.28e-6 NRD=1.16667 NRS=1.16667 M=1
mpm8_3__rcx n45__vdd n36__rst n54__net4 n16__vdd g45p1svt L=45e-9 W=480e-9 AD=76.8e-15 AS=76.8e-15 PD=1.28e-6 PS=1.28e-6 NRD=1.16667 NRS=1.16667 M=1
mpm8_2__rcx n57__net4 n34__rst n45__vdd n16__vdd g45p1svt L=45e-9 W=480e-9 AD=76.8e-15 AS=76.8e-15 PD=1.28e-6 PS=1.28e-6 NRD=1.16667 NRS=1.16667 M=1
mpm8_1__rcx n44__vdd n33__rst n57__net4 n16__vdd g45p1svt L=45e-9 W=480e-9 AD=67.2e-15 AS=67.2e-15 PD=1.26e-6 PS=1.26e-6 NRD=1.16667 NRS=1.16667 M=1
mpm8 n51__net4 n32__rst n52__vdd n16__vdd g45p1svt L=45e-9 W=480e-9 AD=76.8e-15 AS=76.8e-15 PD=1.26e-6 PS=1.26e-6 NRD=1.16667 NRS=1.16667 M=1
mpm3_5__rcx n29__vdd n23__net11 n89__net10 n16__vdd g45p1svt L=45e-9 W=480e-9 AD=76.8e-15 AS=76.8e-15 PD=1.28e-6 PS=1.28e-6 NRD=1.16667 NRS=1.16667 M=1
mpm3_4__rcx n92__net10 n21__net11 n29__vdd n16__vdd g45p1svt L=45e-9 W=480e-9 AD=76.8e-15 AS=76.8e-15 PD=1.28e-6 PS=1.28e-6 NRD=1.16667 NRS=1.16667 M=1
mpm3_3__rcx n27__vdd n19__net11 n92__net10 n16__vdd g45p1svt L=45e-9 W=480e-9 AD=76.8e-15 AS=76.8e-15 PD=1.28e-6 PS=1.28e-6 NRD=1.16667 NRS=1.16667 M=1
mpm3_2__rcx n95__net10 n17__net11 n27__vdd n16__vdd g45p1svt L=45e-9 W=480e-9 AD=76.8e-15 AS=76.8e-15 PD=1.28e-6 PS=1.28e-6 NRD=1.16667 NRS=1.16667 M=1
mpm3_1__rcx n26__vdd n5__net11 n95__net10 n16__vdd g45p1svt L=45e-9 W=480e-9 AD=67.2e-15 AS=67.2e-15 PD=1.26e-6 PS=1.26e-6 NRD=1.16667 NRS=1.16667 M=1
mpm3 n89__net10 n24__net11 n31__vdd n16__vdd g45p1svt L=45e-9 W=480e-9 AD=76.8e-15 AS=76.8e-15 PD=1.26e-6 PS=1.26e-6 NRD=1.16667 NRS=1.16667 M=1
mpm7_5__rcx n37__vdd n47__net4 n49__net3 n16__vdd g45p1svt L=45e-9 W=480e-9 AD=76.8e-15 AS=76.8e-15 PD=1.28e-6 PS=1.28e-6 NRD=1.16667 NRS=1.16667 M=1
mpm7_4__rcx n52__net3 n45__net4 n37__vdd n16__vdd g45p1svt L=45e-9 W=480e-9 AD=76.8e-15 AS=76.8e-15 PD=1.28e-6 PS=1.28e-6 NRD=1.16667 NRS=1.16667 M=1
mpm7_3__rcx n35__vdd n43__net4 n52__net3 n16__vdd g45p1svt L=45e-9 W=480e-9 AD=76.8e-15 AS=76.8e-15 PD=1.28e-6 PS=1.28e-6 NRD=1.16667 NRS=1.16667 M=1
mpm7_2__rcx n55__net3 n41__net4 n35__vdd n16__vdd g45p1svt L=45e-9 W=480e-9 AD=76.8e-15 AS=76.8e-15 PD=1.28e-6 PS=1.28e-6 NRD=1.16667 NRS=1.16667 M=1
mpm7_1__rcx n33__vdd n29__net4 n55__net3 n16__vdd g45p1svt L=45e-9 W=480e-9 AD=67.2e-15 AS=67.2e-15 PD=1.26e-6 PS=1.26e-6 NRD=1.16667 NRS=1.16667 M=1
mpm7 n49__net3 n48__net4 n38__vdd n16__vdd g45p1svt L=45e-9 W=480e-9 AD=76.8e-15 AS=76.8e-15 PD=1.26e-6 PS=1.26e-6 NRD=1.16667 NRS=1.16667 M=1
mi0__i2__pm0 n12__i0__i2__net1 n5__clk n7__i0__net1 n16__vdd g45p1svt L=45e-9 W=120e-9 AD=16.8e-15 AS=16.8e-15 PD=520e-9 PS=520e-9 NRD=1.16667 NRS=1.16667 M=1
mi0__i2__pm2 n92__vdd n2__i0__i2__net2 n9__i0__i2__net1 n16__vdd g45p1svt L=180e-9 W=120e-9 AD=16.8e-15 AS=16.8e-15 PD=520e-9 PS=520e-9 NRD=1.16667 NRS=1.16667 M=1
mi0__i2__pm1_1__rcx n9__i0__i2__net2 n6__i0__i2__net1 n88__vdd n16__vdd g45p1svt L=45e-9 W=480e-9 AD=76.8e-15 AS=76.8e-15 PD=1.26e-6 PS=1.26e-6 NRD=1.16667 NRS=1.16667 M=1
mi0__i2__pm1 n85__vdd n5__i0__i2__net1 n9__i0__i2__net2 n16__vdd g45p1svt L=45e-9 W=480e-9 AD=67.2e-15 AS=67.2e-15 PD=1.26e-6 PS=1.26e-6 NRD=1.16667 NRS=1.16667 M=1
mi0__i2__pm8 n12__i0__i2__net5 n4__i0__net3 n11__i0__i2__net2 n16__vdd g45p1svt L=45e-9 W=120e-9 AD=16.8e-15 AS=16.8e-15 PD=520e-9 PS=520e-9 NRD=1.16667 NRS=1.16667 M=1
mi0__i2__pm10 n82__vdd n2__i0__i2__net4 n9__i0__i2__net5 n16__vdd g45p1svt L=180e-9 W=120e-9 AD=16.8e-15 AS=16.8e-15 PD=520e-9 PS=520e-9 NRD=1.16667 NRS=1.16667 M=1
mi0__i2__pm15 n15__i0__i2__net5 i0__net6 n78__vdd n16__vdd g45p1svt L=45e-9 W=120e-9 AD=16.8e-15 AS=16.8e-15 PD=520e-9 PS=520e-9 NRD=1.16667 NRS=1.16667 M=1
mi0__i2__pm9_1__rcx n10__i0__i2__net4 n6__i0__i2__net5 n75__vdd n16__vdd g45p1svt L=45e-9 W=480e-9 AD=76.8e-15 AS=76.8e-15 PD=1.26e-6 PS=1.26e-6 NRD=1.16667 NRS=1.16667 M=1
mi0__i2__pm9 n72__vdd n5__i0__i2__net5 n10__i0__i2__net4 n16__vdd g45p1svt L=45e-9 W=480e-9 AD=67.2e-15 AS=67.2e-15 PD=1.26e-6 PS=1.26e-6 NRD=1.16667 NRS=1.16667 M=1
mi0__i2__pm11 n28__i0__net1 n6__i0__i2__net4 n69__vdd n16__vdd g45p1svt L=45e-9 W=480e-9 AD=67.2e-15 AS=67.2e-15 PD=1.24e-6 PS=1.24e-6 NRD=1.16667 NRS=1.16667 M=1
mi0__i2__pm13 n19__i0__net7 n17__i0__net1 n66__vdd n16__vdd g45p1svt L=45e-9 W=480e-9 AD=67.2e-15 AS=67.2e-15 PD=1.24e-6 PS=1.24e-6 NRD=1.16667 NRS=1.16667 M=1
mi0__i3__pm0 n13__i0__i3__net1 n2__i0__net7 i0__net8 n16__vdd g45p1svt L=45e-9 W=120e-9 AD=16.8e-15 AS=16.8e-15 PD=520e-9 PS=520e-9 NRD=1.16667 NRS=1.16667 M=1
mi0__i3__pm2 n87__vdd n3__i0__i3__net2 n9__i0__i3__net1 n16__vdd g45p1svt L=180e-9 W=120e-9 AD=16.8e-15 AS=16.8e-15 PD=520e-9 PS=520e-9 NRD=1.16667 NRS=1.16667 M=1
mi0__i3__pm1_1__rcx n11__i0__i3__net2 n7__i0__i3__net1 n84__vdd n16__vdd g45p1svt L=45e-9 W=480e-9 AD=76.8e-15 AS=76.8e-15 PD=1.26e-6 PS=1.26e-6 NRD=1.16667 NRS=1.16667 M=1
mi0__i3__pm1 n81__vdd i0__i3__net1 n11__i0__i3__net2 n16__vdd g45p1svt L=45e-9 W=480e-9 AD=67.2e-15 AS=67.2e-15 PD=1.26e-6 PS=1.26e-6 NRD=1.16667 NRS=1.16667 M=1
mi0__i3__pm8 n13__i0__i3__net5 n4__i0__net1 n6__i0__i3__net2 n16__vdd g45p1svt L=45e-9 W=120e-9 AD=16.8e-15 AS=16.8e-15 PD=520e-9 PS=520e-9 NRD=1.16667 NRS=1.16667 M=1
mi0__i3__pm10 n77__vdd n3__i0__i3__net4 n9__i0__i3__net5 n16__vdd g45p1svt L=180e-9 W=120e-9 AD=16.8e-15 AS=16.8e-15 PD=520e-9 PS=520e-9 NRD=1.16667 NRS=1.16667 M=1
mi0__i3__pm15 n15__i0__i3__net5 n3__i0__net6 n74__vdd n16__vdd g45p1svt L=45e-9 W=120e-9 AD=16.8e-15 AS=16.8e-15 PD=520e-9 PS=520e-9 NRD=1.16667 NRS=1.16667 M=1
mi0__i3__pm9_1__rcx n10__i0__i3__net4 n7__i0__i3__net5 n71__vdd n16__vdd g45p1svt L=45e-9 W=480e-9 AD=76.8e-15 AS=76.8e-15 PD=1.26e-6 PS=1.26e-6 NRD=1.16667 NRS=1.16667 M=1
mi0__i3__pm9 n68__vdd i0__i3__net5 n10__i0__i3__net4 n16__vdd g45p1svt L=45e-9 W=480e-9 AD=67.2e-15 AS=67.2e-15 PD=1.26e-6 PS=1.26e-6 NRD=1.16667 NRS=1.16667 M=1
mi0__i3__pm11 n22__i0__net8 n4__i0__i3__net4 n65__vdd n16__vdd g45p1svt L=45e-9 W=480e-9 AD=67.2e-15 AS=67.2e-15 PD=1.24e-6 PS=1.24e-6 NRD=1.16667 NRS=1.16667 M=1
mi0__i3__pm13 n10__i0__net11 n6__i0__net8 n62__vdd n16__vdd g45p1svt L=45e-9 W=480e-9 AD=67.2e-15 AS=67.2e-15 PD=1.24e-6 PS=1.24e-6 NRD=1.16667 NRS=1.16667 M=1
mi0__i4__pm3 n8__i0__net9 n10__i0__net8 n110__vss n16__vdd g45p1svt L=45e-9 W=240e-9 AD=38.4e-15 AS=38.4e-15 PD=780e-9 PS=780e-9 NRD=1.16667 NRS=1.16667 M=1
mi0__i4__pm2 n55__vdd n2__i0__net11 n8__i0__net9 n16__vdd g45p1svt L=45e-9 W=240e-9 AD=33.6e-15 AS=33.6e-15 PD=780e-9 PS=780e-9 NRD=1.16667 NRS=1.16667 M=1
mi0__i4__pm6 n9__i0__net10 n5__i0__net9 n50__vdd n16__vdd g45p1svt L=45e-9 W=480e-9 AD=67.2e-15 AS=67.2e-15 PD=1.24e-6 PS=1.24e-6 NRD=1.16667 NRS=1.16667 M=1
mi0__i4__pm5 n47__vdd n5__i0__net10 n16__i0__net9 n16__vdd g45p1svt L=45e-9 W=480e-9 AD=67.2e-15 AS=67.2e-15 PD=1.24e-6 PS=1.24e-6 NRD=1.16667 NRS=1.16667 M=1
mi0__i4__pm0 n16__i0__net10 n15__i0__net8 n41__vdd n16__vdd g45p1svt L=45e-9 W=240e-9 AD=38.4e-15 AS=38.4e-15 PD=780e-9 PS=780e-9 NRD=1.16667 NRS=1.16667 M=1
mi0__i4__pm1 n130__vss n6__i0__net11 n16__i0__net10 n16__vdd g45p1svt L=45e-9 W=240e-9 AD=33.6e-15 AS=33.6e-15 PD=780e-9 PS=780e-9 NRD=1.16667 NRS=1.16667 M=1
mi0__pm17 n25__net7 n4__i0__net9 n58__vdd n16__vdd g45p1svt L=45e-9 W=480e-9 AD=67.2e-15 AS=67.2e-15 PD=1.24e-6 PS=1.24e-6 NRD=1.16667 NRS=1.16667 M=1
mi0__pm16 n26__net11 n4__i0__net10 n63__vdd n16__vdd g45p1svt L=45e-9 W=480e-9 AD=67.2e-15 AS=67.2e-15 PD=1.24e-6 PS=1.24e-6 NRD=1.16667 NRS=1.16667 M=1
mi0__pm1 n5__i0__net6 n1__rst n91__vdd n16__vdd g45p1svt L=45e-9 W=240e-9 AD=33.6e-15 AS=33.6e-15 PD=760e-9 PS=760e-9 NRD=1.16667 NRS=1.16667 M=1
mi0__pm0 n7__i0__net3 n3__clk n93__vdd n16__vdd g45p1svt L=45e-9 W=240e-9 AD=33.6e-15 AS=33.6e-15 PD=760e-9 PS=760e-9 NRD=1.16667 NRS=1.16667 M=1
mi7__pm0 n12__i7__net1 n42__net10 n5__y_in_3 n97__vdd g45p1svt L=45e-9 W=120e-9 AD=16.8e-15 AS=16.8e-15 PD=520e-9 PS=520e-9 NRD=1.16667 NRS=1.16667 M=1
mi7__pm2 n130__vdd n2__i7__net2 n9__i7__net1 n97__vdd g45p1svt L=180e-9 W=120e-9 AD=16.8e-15 AS=16.8e-15 PD=520e-9 PS=520e-9 NRD=1.16667 NRS=1.16667 M=1
mi7__pm1_1__rcx n8__i7__net2 n6__i7__net1 n128__vdd n97__vdd g45p1svt L=45e-9 W=480e-9 AD=76.8e-15 AS=76.8e-15 PD=1.26e-6 PS=1.26e-6 NRD=1.16667 NRS=1.16667 M=1
mi7__pm1 n126__vdd n5__i7__net1 n8__i7__net2 n97__vdd g45p1svt L=45e-9 W=480e-9 AD=67.2e-15 AS=67.2e-15 PD=1.26e-6 PS=1.26e-6 NRD=1.16667 NRS=1.16667 M=1
mi7__pm8 n12__i7__net5 n50__net9 n10__i7__net2 n97__vdd g45p1svt L=45e-9 W=120e-9 AD=16.8e-15 AS=16.8e-15 PD=520e-9 PS=520e-9 NRD=1.16667 NRS=1.16667 M=1
mi7__pm10 n124__vdd n2__i7__net4 n9__i7__net5 n97__vdd g45p1svt L=180e-9 W=120e-9 AD=16.8e-15 AS=16.8e-15 PD=520e-9 PS=520e-9 NRD=1.16667 NRS=1.16667 M=1
mi7__pm15 n15__i7__net5 n21__net4 n122__vdd n97__vdd g45p1svt L=45e-9 W=120e-9 AD=16.8e-15 AS=16.8e-15 PD=520e-9 PS=520e-9 NRD=1.16667 NRS=1.16667 M=1
mi7__pm9_1__rcx n10__i7__net4 n6__i7__net5 n120__vdd n97__vdd g45p1svt L=45e-9 W=480e-9 AD=76.8e-15 AS=76.8e-15 PD=1.26e-6 PS=1.26e-6 NRD=1.16667 NRS=1.16667 M=1
mi7__pm9 n118__vdd n5__i7__net5 n10__i7__net4 n97__vdd g45p1svt L=45e-9 W=480e-9 AD=67.2e-15 AS=67.2e-15 PD=1.26e-6 PS=1.26e-6 NRD=1.16667 NRS=1.16667 M=1
mi7__pm11 n7__y_out_b_3 n6__i7__net4 n116__vdd n97__vdd g45p1svt L=45e-9 W=480e-9 AD=67.2e-15 AS=67.2e-15 PD=1.24e-6 PS=1.24e-6 NRD=1.16667 NRS=1.16667 M=1
mi7__pm13 n3__y_out_3 n4__y_out_b_3 n94__vdd n97__vdd g45p1svt L=45e-9 W=480e-9 AD=67.2e-15 AS=67.2e-15 PD=1.24e-6 PS=1.24e-6 NRD=1.16667 NRS=1.16667 M=1
mi1__pm0 n12__i1__net1 n2__net10 n3__x_in_3 n97__vdd g45p1svt L=45e-9 W=120e-9 AD=16.8e-15 AS=16.8e-15 PD=520e-9 PS=520e-9 NRD=1.16667 NRS=1.16667 M=1
mi1__pm2 n153__vdd n2__i1__net2 n9__i1__net1 n97__vdd g45p1svt L=180e-9 W=120e-9 AD=16.8e-15 AS=16.8e-15 PD=520e-9 PS=520e-9 NRD=1.16667 NRS=1.16667 M=1
mi1__pm1_1__rcx n9__i1__net2 n6__i1__net1 n151__vdd n97__vdd g45p1svt L=45e-9 W=480e-9 AD=76.8e-15 AS=76.8e-15 PD=1.26e-6 PS=1.26e-6 NRD=1.16667 NRS=1.16667 M=1
mi1__pm1 n147__vdd n5__i1__net1 n9__i1__net2 n97__vdd g45p1svt L=45e-9 W=480e-9 AD=67.2e-15 AS=67.2e-15 PD=1.26e-6 PS=1.26e-6 NRD=1.16667 NRS=1.16667 M=1
mi1__pm8 n12__i1__net5 n10__net9 n11__i1__net2 n97__vdd g45p1svt L=45e-9 W=120e-9 AD=16.8e-15 AS=16.8e-15 PD=520e-9 PS=520e-9 NRD=1.16667 NRS=1.16667 M=1
mi1__pm10 n144__vdd n2__i1__net4 n9__i1__net5 n97__vdd g45p1svt L=180e-9 W=120e-9 AD=16.8e-15 AS=16.8e-15 PD=520e-9 PS=520e-9 NRD=1.16667 NRS=1.16667 M=1
mi1__pm15 n15__i1__net5 net4 n140__vdd n97__vdd g45p1svt L=45e-9 W=120e-9 AD=16.8e-15 AS=16.8e-15 PD=520e-9 PS=520e-9 NRD=1.16667 NRS=1.16667 M=1
mi1__pm9_1__rcx n10__i1__net4 n6__i1__net5 n138__vdd n97__vdd g45p1svt L=45e-9 W=480e-9 AD=76.8e-15 AS=76.8e-15 PD=1.26e-6 PS=1.26e-6 NRD=1.16667 NRS=1.16667 M=1
mi1__pm9 n136__vdd n5__i1__net5 n10__i1__net4 n97__vdd g45p1svt L=45e-9 W=480e-9 AD=67.2e-15 AS=67.2e-15 PD=1.26e-6 PS=1.26e-6 NRD=1.16667 NRS=1.16667 M=1
mi1__pm11 n7__x_out_b_3 n6__i1__net4 n134__vdd n97__vdd g45p1svt L=45e-9 W=480e-9 AD=67.2e-15 AS=67.2e-15 PD=1.24e-6 PS=1.24e-6 NRD=1.16667 NRS=1.16667 M=1
mi1__pm13 n3__x_out_3 n4__x_out_b_3 n132__vdd n97__vdd g45p1svt L=45e-9 W=480e-9 AD=67.2e-15 AS=67.2e-15 PD=1.24e-6 PS=1.24e-6 NRD=1.16667 NRS=1.16667 M=1
mi4__pm0 n12__i4__net1 n46__net10 n5__y_in_1 n157__vdd g45p1svt L=45e-9 W=120e-9 AD=16.8e-15 AS=16.8e-15 PD=520e-9 PS=520e-9 NRD=1.16667 NRS=1.16667 M=1
mi4__pm2 n190__vdd n2__i4__net2 n9__i4__net1 n157__vdd g45p1svt L=180e-9 W=120e-9 AD=16.8e-15 AS=16.8e-15 PD=520e-9 PS=520e-9 NRD=1.16667 NRS=1.16667 M=1
mi4__pm1_1__rcx n8__i4__net2 n6__i4__net1 n188__vdd n157__vdd g45p1svt L=45e-9 W=480e-9 AD=76.8e-15 AS=76.8e-15 PD=1.26e-6 PS=1.26e-6 NRD=1.16667 NRS=1.16667 M=1
mi4__pm1 n186__vdd n5__i4__net1 n8__i4__net2 n157__vdd g45p1svt L=45e-9 W=480e-9 AD=67.2e-15 AS=67.2e-15 PD=1.26e-6 PS=1.26e-6 NRD=1.16667 NRS=1.16667 M=1
mi4__pm8 n12__i4__net5 n54__net9 n10__i4__net2 n157__vdd g45p1svt L=45e-9 W=120e-9 AD=16.8e-15 AS=16.8e-15 PD=520e-9 PS=520e-9 NRD=1.16667 NRS=1.16667 M=1
mi4__pm10 n184__vdd n2__i4__net4 n9__i4__net5 n157__vdd g45p1svt L=180e-9 W=120e-9 AD=16.8e-15 AS=16.8e-15 PD=520e-9 PS=520e-9 NRD=1.16667 NRS=1.16667 M=1
mi4__pm15 n15__i4__net5 n25__net4 n182__vdd n157__vdd g45p1svt L=45e-9 W=120e-9 AD=16.8e-15 AS=16.8e-15 PD=520e-9 PS=520e-9 NRD=1.16667 NRS=1.16667 M=1
mi4__pm9_1__rcx n10__i4__net4 n6__i4__net5 n180__vdd n157__vdd g45p1svt L=45e-9 W=480e-9 AD=76.8e-15 AS=76.8e-15 PD=1.26e-6 PS=1.26e-6 NRD=1.16667 NRS=1.16667 M=1
mi4__pm9 n178__vdd n5__i4__net5 n10__i4__net4 n157__vdd g45p1svt L=45e-9 W=480e-9 AD=67.2e-15 AS=67.2e-15 PD=1.26e-6 PS=1.26e-6 NRD=1.16667 NRS=1.16667 M=1
mi4__pm11 n7__y_out_b_1 n6__i4__net4 n176__vdd n157__vdd g45p1svt L=45e-9 W=480e-9 AD=67.2e-15 AS=67.2e-15 PD=1.24e-6 PS=1.24e-6 NRD=1.16667 NRS=1.16667 M=1
mi4__pm13 n3__y_out_1 n4__y_out_b_1 n154__vdd n157__vdd g45p1svt L=45e-9 W=480e-9 AD=67.2e-15 AS=67.2e-15 PD=1.24e-6 PS=1.24e-6 NRD=1.16667 NRS=1.16667 M=1
mi3__pm0 n12__i3__net1 n6__net10 n3__x_in_1 n157__vdd g45p1svt L=45e-9 W=120e-9 AD=16.8e-15 AS=16.8e-15 PD=520e-9 PS=520e-9 NRD=1.16667 NRS=1.16667 M=1
mi3__pm2 n213__vdd n2__i3__net2 n9__i3__net1 n157__vdd g45p1svt L=180e-9 W=120e-9 AD=16.8e-15 AS=16.8e-15 PD=520e-9 PS=520e-9 NRD=1.16667 NRS=1.16667 M=1
mi3__pm1_1__rcx n9__i3__net2 n6__i3__net1 n211__vdd n157__vdd g45p1svt L=45e-9 W=480e-9 AD=76.8e-15 AS=76.8e-15 PD=1.26e-6 PS=1.26e-6 NRD=1.16667 NRS=1.16667 M=1
mi3__pm1 n207__vdd n5__i3__net1 n9__i3__net2 n157__vdd g45p1svt L=45e-9 W=480e-9 AD=67.2e-15 AS=67.2e-15 PD=1.26e-6 PS=1.26e-6 NRD=1.16667 NRS=1.16667 M=1
mi3__pm8 n12__i3__net5 n14__net9 n11__i3__net2 n157__vdd g45p1svt L=45e-9 W=120e-9 AD=16.8e-15 AS=16.8e-15 PD=520e-9 PS=520e-9 NRD=1.16667 NRS=1.16667 M=1
mi3__pm10 n204__vdd n2__i3__net4 n9__i3__net5 n157__vdd g45p1svt L=180e-9 W=120e-9 AD=16.8e-15 AS=16.8e-15 PD=520e-9 PS=520e-9 NRD=1.16667 NRS=1.16667 M=1
mi3__pm15 n15__i3__net5 n5__net4 n200__vdd n157__vdd g45p1svt L=45e-9 W=120e-9 AD=16.8e-15 AS=16.8e-15 PD=520e-9 PS=520e-9 NRD=1.16667 NRS=1.16667 M=1
mi3__pm9_1__rcx n10__i3__net4 n6__i3__net5 n198__vdd n157__vdd g45p1svt L=45e-9 W=480e-9 AD=76.8e-15 AS=76.8e-15 PD=1.26e-6 PS=1.26e-6 NRD=1.16667 NRS=1.16667 M=1
mi3__pm9 n196__vdd n5__i3__net5 n10__i3__net4 n157__vdd g45p1svt L=45e-9 W=480e-9 AD=67.2e-15 AS=67.2e-15 PD=1.26e-6 PS=1.26e-6 NRD=1.16667 NRS=1.16667 M=1
mi3__pm11 n7__x_out_b_1 n6__i3__net4 n194__vdd n157__vdd g45p1svt L=45e-9 W=480e-9 AD=67.2e-15 AS=67.2e-15 PD=1.24e-6 PS=1.24e-6 NRD=1.16667 NRS=1.16667 M=1
mi3__pm13 n3__x_out_1 n4__x_out_b_1 n192__vdd n157__vdd g45p1svt L=45e-9 W=480e-9 AD=67.2e-15 AS=67.2e-15 PD=1.24e-6 PS=1.24e-6 NRD=1.16667 NRS=1.16667 M=1
mi6__pm0 n13__i6__net1 n44__net10 n3__y_in_2 n97__vdd g45p1svt L=45e-9 W=120e-9 AD=16.8e-15 AS=16.8e-15 PD=520e-9 PS=520e-9 NRD=1.16667 NRS=1.16667 M=1
mi6__pm2 n129__vdd n3__i6__net2 n9__i6__net1 n97__vdd g45p1svt L=180e-9 W=120e-9 AD=16.8e-15 AS=16.8e-15 PD=520e-9 PS=520e-9 NRD=1.16667 NRS=1.16667 M=1
mi6__pm1_1__rcx n10__i6__net2 n7__i6__net1 n127__vdd n97__vdd g45p1svt L=45e-9 W=480e-9 AD=76.8e-15 AS=76.8e-15 PD=1.26e-6 PS=1.26e-6 NRD=1.16667 NRS=1.16667 M=1
mi6__pm1 n125__vdd i6__net1 n10__i6__net2 n97__vdd g45p1svt L=45e-9 W=480e-9 AD=67.2e-15 AS=67.2e-15 PD=1.26e-6 PS=1.26e-6 NRD=1.16667 NRS=1.16667 M=1
mi6__pm8 n13__i6__net5 n52__net9 n5__i6__net2 n97__vdd g45p1svt L=45e-9 W=120e-9 AD=16.8e-15 AS=16.8e-15 PD=520e-9 PS=520e-9 NRD=1.16667 NRS=1.16667 M=1
mi6__pm10 n123__vdd n3__i6__net4 n9__i6__net5 n97__vdd g45p1svt L=180e-9 W=120e-9 AD=16.8e-15 AS=16.8e-15 PD=520e-9 PS=520e-9 NRD=1.16667 NRS=1.16667 M=1
mi6__pm15 n15__i6__net5 n23__net4 n121__vdd n97__vdd g45p1svt L=45e-9 W=120e-9 AD=16.8e-15 AS=16.8e-15 PD=520e-9 PS=520e-9 NRD=1.16667 NRS=1.16667 M=1
mi6__pm9_1__rcx n10__i6__net4 n7__i6__net5 n119__vdd n97__vdd g45p1svt L=45e-9 W=480e-9 AD=76.8e-15 AS=76.8e-15 PD=1.26e-6 PS=1.26e-6 NRD=1.16667 NRS=1.16667 M=1
mi6__pm9 n117__vdd i6__net5 n10__i6__net4 n97__vdd g45p1svt L=45e-9 W=480e-9 AD=67.2e-15 AS=67.2e-15 PD=1.26e-6 PS=1.26e-6 NRD=1.16667 NRS=1.16667 M=1
mi6__pm11 n8__y_out_b_2 n4__i6__net4 n115__vdd n97__vdd g45p1svt L=45e-9 W=480e-9 AD=67.2e-15 AS=67.2e-15 PD=1.24e-6 PS=1.24e-6 NRD=1.16667 NRS=1.16667 M=1
mi6__pm13 n1__y_out_2 n1__y_out_b_2 n114__vdd n97__vdd g45p1svt L=45e-9 W=480e-9 AD=67.2e-15 AS=67.2e-15 PD=1.24e-6 PS=1.24e-6 NRD=1.16667 NRS=1.16667 M=1
mi2__pm0 n13__i2__net1 n4__net10 n1__x_in_2 n97__vdd g45p1svt L=45e-9 W=120e-9 AD=16.8e-15 AS=16.8e-15 PD=520e-9 PS=520e-9 NRD=1.16667 NRS=1.16667 M=1
mi2__pm2 n150__vdd n3__i2__net2 n9__i2__net1 n97__vdd g45p1svt L=180e-9 W=120e-9 AD=16.8e-15 AS=16.8e-15 PD=520e-9 PS=520e-9 NRD=1.16667 NRS=1.16667 M=1
mi2__pm1_1__rcx n11__i2__net2 n7__i2__net1 n146__vdd n97__vdd g45p1svt L=45e-9 W=480e-9 AD=76.8e-15 AS=76.8e-15 PD=1.26e-6 PS=1.26e-6 NRD=1.16667 NRS=1.16667 M=1
mi2__pm1 n143__vdd i2__net1 n11__i2__net2 n97__vdd g45p1svt L=45e-9 W=480e-9 AD=67.2e-15 AS=67.2e-15 PD=1.26e-6 PS=1.26e-6 NRD=1.16667 NRS=1.16667 M=1
mi2__pm8 n13__i2__net5 n12__net9 n6__i2__net2 n97__vdd g45p1svt L=45e-9 W=120e-9 AD=16.8e-15 AS=16.8e-15 PD=520e-9 PS=520e-9 NRD=1.16667 NRS=1.16667 M=1
mi2__pm10 n141__vdd n3__i2__net4 n9__i2__net5 n97__vdd g45p1svt L=180e-9 W=120e-9 AD=16.8e-15 AS=16.8e-15 PD=520e-9 PS=520e-9 NRD=1.16667 NRS=1.16667 M=1
mi2__pm15 n15__i2__net5 n3__net4 n139__vdd n97__vdd g45p1svt L=45e-9 W=120e-9 AD=16.8e-15 AS=16.8e-15 PD=520e-9 PS=520e-9 NRD=1.16667 NRS=1.16667 M=1
mi2__pm9_1__rcx n10__i2__net4 n7__i2__net5 n137__vdd n97__vdd g45p1svt L=45e-9 W=480e-9 AD=76.8e-15 AS=76.8e-15 PD=1.26e-6 PS=1.26e-6 NRD=1.16667 NRS=1.16667 M=1
mi2__pm9 n135__vdd i2__net5 n10__i2__net4 n97__vdd g45p1svt L=45e-9 W=480e-9 AD=67.2e-15 AS=67.2e-15 PD=1.26e-6 PS=1.26e-6 NRD=1.16667 NRS=1.16667 M=1
mi2__pm11 n8__x_out_b_2 n4__i2__net4 n133__vdd n97__vdd g45p1svt L=45e-9 W=480e-9 AD=67.2e-15 AS=67.2e-15 PD=1.24e-6 PS=1.24e-6 NRD=1.16667 NRS=1.16667 M=1
mi2__pm13 n1__x_out_2 n1__x_out_b_2 n131__vdd n97__vdd g45p1svt L=45e-9 W=480e-9 AD=67.2e-15 AS=67.2e-15 PD=1.24e-6 PS=1.24e-6 NRD=1.16667 NRS=1.16667 M=1
mi5__pm0 n13__i5__net1 n48__net10 n3__y_in_0 n157__vdd g45p1svt L=45e-9 W=120e-9 AD=16.8e-15 AS=16.8e-15 PD=520e-9 PS=520e-9 NRD=1.16667 NRS=1.16667 M=1
mi5__pm2 n189__vdd n3__i5__net2 n9__i5__net1 n157__vdd g45p1svt L=180e-9 W=120e-9 AD=16.8e-15 AS=16.8e-15 PD=520e-9 PS=520e-9 NRD=1.16667 NRS=1.16667 M=1
mi5__pm1_1__rcx n10__i5__net2 n7__i5__net1 n187__vdd n157__vdd g45p1svt L=45e-9 W=480e-9 AD=76.8e-15 AS=76.8e-15 PD=1.26e-6 PS=1.26e-6 NRD=1.16667 NRS=1.16667 M=1
mi5__pm1 n185__vdd i5__net1 n10__i5__net2 n157__vdd g45p1svt L=45e-9 W=480e-9 AD=67.2e-15 AS=67.2e-15 PD=1.26e-6 PS=1.26e-6 NRD=1.16667 NRS=1.16667 M=1
mi5__pm8 n13__i5__net5 n56__net9 n5__i5__net2 n157__vdd g45p1svt L=45e-9 W=120e-9 AD=16.8e-15 AS=16.8e-15 PD=520e-9 PS=520e-9 NRD=1.16667 NRS=1.16667 M=1
mi5__pm10 n183__vdd n3__i5__net4 n9__i5__net5 n157__vdd g45p1svt L=180e-9 W=120e-9 AD=16.8e-15 AS=16.8e-15 PD=520e-9 PS=520e-9 NRD=1.16667 NRS=1.16667 M=1
mi5__pm15 n15__i5__net5 n27__net4 n181__vdd n157__vdd g45p1svt L=45e-9 W=120e-9 AD=16.8e-15 AS=16.8e-15 PD=520e-9 PS=520e-9 NRD=1.16667 NRS=1.16667 M=1
mi5__pm9_1__rcx n10__i5__net4 n7__i5__net5 n179__vdd n157__vdd g45p1svt L=45e-9 W=480e-9 AD=76.8e-15 AS=76.8e-15 PD=1.26e-6 PS=1.26e-6 NRD=1.16667 NRS=1.16667 M=1
mi5__pm9 n177__vdd i5__net5 n10__i5__net4 n157__vdd g45p1svt L=45e-9 W=480e-9 AD=67.2e-15 AS=67.2e-15 PD=1.26e-6 PS=1.26e-6 NRD=1.16667 NRS=1.16667 M=1
mi5__pm11 n8__y_out_b_0 n4__i5__net4 n175__vdd n157__vdd g45p1svt L=45e-9 W=480e-9 AD=67.2e-15 AS=67.2e-15 PD=1.24e-6 PS=1.24e-6 NRD=1.16667 NRS=1.16667 M=1
mi5__pm13 n1__y_out_0 n1__y_out_b_0 n174__vdd n157__vdd g45p1svt L=45e-9 W=480e-9 AD=67.2e-15 AS=67.2e-15 PD=1.24e-6 PS=1.24e-6 NRD=1.16667 NRS=1.16667 M=1
mi8__pm0 n13__i8__net1 n8__net10 n1__x_in_0 n157__vdd g45p1svt L=45e-9 W=120e-9 AD=16.8e-15 AS=16.8e-15 PD=520e-9 PS=520e-9 NRD=1.16667 NRS=1.16667 M=1
mi8__pm2 n210__vdd n3__i8__net2 n9__i8__net1 n157__vdd g45p1svt L=180e-9 W=120e-9 AD=16.8e-15 AS=16.8e-15 PD=520e-9 PS=520e-9 NRD=1.16667 NRS=1.16667 M=1
mi8__pm1_1__rcx n11__i8__net2 n7__i8__net1 n206__vdd n157__vdd g45p1svt L=45e-9 W=480e-9 AD=76.8e-15 AS=76.8e-15 PD=1.26e-6 PS=1.26e-6 NRD=1.16667 NRS=1.16667 M=1
mi8__pm1 n203__vdd i8__net1 n11__i8__net2 n157__vdd g45p1svt L=45e-9 W=480e-9 AD=67.2e-15 AS=67.2e-15 PD=1.26e-6 PS=1.26e-6 NRD=1.16667 NRS=1.16667 M=1
mi8__pm8 n13__i8__net5 n16__net9 n6__i8__net2 n157__vdd g45p1svt L=45e-9 W=120e-9 AD=16.8e-15 AS=16.8e-15 PD=520e-9 PS=520e-9 NRD=1.16667 NRS=1.16667 M=1
mi8__pm10 n201__vdd n3__i8__net4 n9__i8__net5 n157__vdd g45p1svt L=180e-9 W=120e-9 AD=16.8e-15 AS=16.8e-15 PD=520e-9 PS=520e-9 NRD=1.16667 NRS=1.16667 M=1
mi8__pm15 n15__i8__net5 n7__net4 n199__vdd n157__vdd g45p1svt L=45e-9 W=120e-9 AD=16.8e-15 AS=16.8e-15 PD=520e-9 PS=520e-9 NRD=1.16667 NRS=1.16667 M=1
mi8__pm9_1__rcx n10__i8__net4 n7__i8__net5 n197__vdd n157__vdd g45p1svt L=45e-9 W=480e-9 AD=76.8e-15 AS=76.8e-15 PD=1.26e-6 PS=1.26e-6 NRD=1.16667 NRS=1.16667 M=1
mi8__pm9 n195__vdd i8__net5 n10__i8__net4 n157__vdd g45p1svt L=45e-9 W=480e-9 AD=67.2e-15 AS=67.2e-15 PD=1.26e-6 PS=1.26e-6 NRD=1.16667 NRS=1.16667 M=1
mi8__pm11 n8__x_out_b_0 n4__i8__net4 n193__vdd n157__vdd g45p1svt L=45e-9 W=480e-9 AD=67.2e-15 AS=67.2e-15 PD=1.24e-6 PS=1.24e-6 NRD=1.16667 NRS=1.16667 M=1
mi8__pm13 n1__x_out_0 n1__x_out_b_0 n191__vdd n157__vdd g45p1svt L=45e-9 W=480e-9 AD=67.2e-15 AS=67.2e-15 PD=1.24e-6 PS=1.24e-6 NRD=1.16667 NRS=1.16667 M=1
mpm9 n2__clk_div4_out n4__net11 n34__vdd n16__vdd g45p1svt L=45e-9 W=480e-9 AD=67.2e-15 AS=67.2e-15 PD=1.24e-6 PS=1.24e-6 NRD=1.16667 NRS=1.16667 M=1
mpm10 n1__clk_div4_out_b n4__net7 n36__vdd n16__vdd g45p1svt L=45e-9 W=480e-9 AD=67.2e-15 AS=67.2e-15 PD=1.24e-6 PS=1.24e-6 NRD=1.16667 NRS=1.16667 M=1
mnm0_5__rcx n10__vss n23__net7 n73__net9 n3__vss g45n1svt L=45e-9 W=240e-9 AD=38.4e-15 AS=38.4e-15 PD=800e-9 PS=800e-9 NRD=1.16667 NRS=1.16667 M=1
mnm0_4__rcx n76__net9 n21__net7 n10__vss n3__vss g45n1svt L=45e-9 W=240e-9 AD=38.4e-15 AS=38.4e-15 PD=800e-9 PS=800e-9 NRD=1.16667 NRS=1.16667 M=1
mnm0_3__rcx n9__vss n19__net7 n76__net9 n3__vss g45n1svt L=45e-9 W=240e-9 AD=38.4e-15 AS=38.4e-15 PD=800e-9 PS=800e-9 NRD=1.16667 NRS=1.16667 M=1
mnm0_2__rcx n79__net9 n17__net7 n9__vss n3__vss g45n1svt L=45e-9 W=240e-9 AD=38.4e-15 AS=38.4e-15 PD=800e-9 PS=800e-9 NRD=1.16667 NRS=1.16667 M=1
mnm0_1__rcx n1__vss n5__net7 n79__net9 n3__vss g45n1svt L=45e-9 W=240e-9 AD=33.6e-15 AS=33.6e-15 PD=780e-9 PS=780e-9 NRD=1.16667 NRS=1.16667 M=1
mnm0 n73__net9 n24__net7 n11__vss n3__vss g45n1svt L=45e-9 W=240e-9 AD=38.4e-15 AS=38.4e-15 PD=780e-9 PS=780e-9 NRD=1.16667 NRS=1.16667 M=1
mnm8_5__rcx n18__vss n41__rst n49__net4 n3__vss g45n1svt L=45e-9 W=240e-9 AD=38.4e-15 AS=38.4e-15 PD=800e-9 PS=800e-9 NRD=1.16667 NRS=1.16667 M=1
mnm8_4__rcx n52__net4 n39__rst n18__vss n3__vss g45n1svt L=45e-9 W=240e-9 AD=38.4e-15 AS=38.4e-15 PD=800e-9 PS=800e-9 NRD=1.16667 NRS=1.16667 M=1
mnm8_3__rcx n16__vss n37__rst n52__net4 n3__vss g45n1svt L=45e-9 W=240e-9 AD=38.4e-15 AS=38.4e-15 PD=800e-9 PS=800e-9 NRD=1.16667 NRS=1.16667 M=1
mnm8_2__rcx n55__net4 n35__rst n16__vss n3__vss g45n1svt L=45e-9 W=240e-9 AD=38.4e-15 AS=38.4e-15 PD=800e-9 PS=800e-9 NRD=1.16667 NRS=1.16667 M=1
mnm8_1__rcx n14__vss n23__rst n55__net4 n3__vss g45n1svt L=45e-9 W=240e-9 AD=33.6e-15 AS=33.6e-15 PD=780e-9 PS=780e-9 NRD=1.16667 NRS=1.16667 M=1
mnm8 n49__net4 n42__rst n20__vss n3__vss g45n1svt L=45e-9 W=240e-9 AD=38.4e-15 AS=38.4e-15 PD=780e-9 PS=780e-9 NRD=1.16667 NRS=1.16667 M=1
mnm1_5__rcx n91__vss n22__net11 n91__net10 n3__vss g45n1svt L=45e-9 W=240e-9 AD=38.4e-15 AS=38.4e-15 PD=800e-9 PS=800e-9 NRD=1.16667 NRS=1.16667 M=1
mnm1_4__rcx n94__net10 n20__net11 n91__vss n3__vss g45n1svt L=45e-9 W=240e-9 AD=38.4e-15 AS=38.4e-15 PD=800e-9 PS=800e-9 NRD=1.16667 NRS=1.16667 M=1
mnm1_3__rcx n89__vss n18__net11 n94__net10 n3__vss g45n1svt L=45e-9 W=240e-9 AD=38.4e-15 AS=38.4e-15 PD=800e-9 PS=800e-9 NRD=1.16667 NRS=1.16667 M=1
mnm1_2__rcx n97__net10 n16__net11 n89__vss n3__vss g45n1svt L=45e-9 W=240e-9 AD=38.4e-15 AS=38.4e-15 PD=800e-9 PS=800e-9 NRD=1.16667 NRS=1.16667 M=1
mnm1_1__rcx n47__vss n15__net11 n97__net10 n3__vss g45n1svt L=45e-9 W=240e-9 AD=33.6e-15 AS=33.6e-15 PD=780e-9 PS=780e-9 NRD=1.16667 NRS=1.16667 M=1
mnm1 n91__net10 n14__net11 n93__vss n3__vss g45n1svt L=45e-9 W=240e-9 AD=38.4e-15 AS=38.4e-15 PD=780e-9 PS=780e-9 NRD=1.16667 NRS=1.16667 M=1
mnm7_5__rcx n98__vss n46__net4 n51__net3 n3__vss g45n1svt L=45e-9 W=240e-9 AD=38.4e-15 AS=38.4e-15 PD=800e-9 PS=800e-9 NRD=1.16667 NRS=1.16667 M=1
mnm7_4__rcx n54__net3 n44__net4 n98__vss n3__vss g45n1svt L=45e-9 W=240e-9 AD=38.4e-15 AS=38.4e-15 PD=800e-9 PS=800e-9 NRD=1.16667 NRS=1.16667 M=1
mnm7_3__rcx n97__vss n42__net4 n54__net3 n3__vss g45n1svt L=45e-9 W=240e-9 AD=38.4e-15 AS=38.4e-15 PD=800e-9 PS=800e-9 NRD=1.16667 NRS=1.16667 M=1
mnm7_2__rcx n57__net3 n40__net4 n97__vss n3__vss g45n1svt L=45e-9 W=240e-9 AD=38.4e-15 AS=38.4e-15 PD=800e-9 PS=800e-9 NRD=1.16667 NRS=1.16667 M=1
mnm7_1__rcx n95__vss n39__net4 n57__net3 n3__vss g45n1svt L=45e-9 W=240e-9 AD=33.6e-15 AS=33.6e-15 PD=780e-9 PS=780e-9 NRD=1.16667 NRS=1.16667 M=1
mnm7 n51__net3 n38__net4 n99__vss n3__vss g45n1svt L=45e-9 W=240e-9 AD=38.4e-15 AS=38.4e-15 PD=780e-9 PS=780e-9 NRD=1.16667 NRS=1.16667 M=1
mi0__i2__nm0 n13__i0__i2__net1 n2__i0__net3 n5__i0__net1 n3__vss g45n1svt L=45e-9 W=120e-9 AD=16.8e-15 AS=16.8e-15 PD=520e-9 PS=520e-9 NRD=1.16667 NRS=1.16667 M=1
mi0__i2__nm8 n44__vss n3__i0__i2__net2 n8__i0__i2__net1 n3__vss g45n1svt L=570e-9 W=120e-9 AD=16.8e-15 AS=16.8e-15 PD=520e-9 PS=520e-9 NRD=1.16667 NRS=1.16667 M=1
mi0__i2__nm18 n42__vss n5__rst n15__i0__i2__net1 n3__vss g45n1svt L=45e-9 W=120e-9 AD=16.8e-15 AS=16.8e-15 PD=520e-9 PS=520e-9 NRD=1.16667 NRS=1.16667 M=1
mi0__i2__nm2_1__rcx n12__i0__i2__net2 n7__i0__i2__net1 n40__vss n3__vss g45n1svt L=45e-9 W=240e-9 AD=38.4e-15 AS=38.4e-15 PD=780e-9 PS=780e-9 NRD=1.16667 NRS=1.16667 M=1
mi0__i2__nm2 n38__vss i0__i2__net1 n12__i0__i2__net2 n3__vss g45n1svt L=45e-9 W=240e-9 AD=33.6e-15 AS=33.6e-15 PD=780e-9 PS=780e-9 NRD=1.16667 NRS=1.16667 M=1
mi0__i2__nm12 n13__i0__i2__net5 n7__clk n6__i0__i2__net2 n3__vss g45n1svt L=45e-9 W=120e-9 AD=16.8e-15 AS=16.8e-15 PD=520e-9 PS=520e-9 NRD=1.16667 NRS=1.16667 M=1
mi0__i2__nm15 n35__vss n3__i0__i2__net4 n8__i0__i2__net5 n3__vss g45n1svt L=570e-9 W=120e-9 AD=16.8e-15 AS=16.8e-15 PD=520e-9 PS=520e-9 NRD=1.16667 NRS=1.16667 M=1
mi0__i2__nm13_1__rcx n8__i0__i2__net4 n7__i0__i2__net5 n33__vss n3__vss g45n1svt L=45e-9 W=240e-9 AD=38.4e-15 AS=38.4e-15 PD=780e-9 PS=780e-9 NRD=1.16667 NRS=1.16667 M=1
mi0__i2__nm13 n31__vss i0__i2__net5 n8__i0__i2__net4 n3__vss g45n1svt L=45e-9 W=240e-9 AD=33.6e-15 AS=33.6e-15 PD=780e-9 PS=780e-9 NRD=1.16667 NRS=1.16667 M=1
mi0__i2__nm16 n29__i0__net1 n4__i0__i2__net4 n29__vss n3__vss g45n1svt L=45e-9 W=240e-9 AD=33.6e-15 AS=33.6e-15 PD=760e-9 PS=760e-9 NRD=1.16667 NRS=1.16667 M=1
mi0__i2__nm17 n17__i0__net7 n14__i0__net1 n27__vss n3__vss g45n1svt L=45e-9 W=240e-9 AD=33.6e-15 AS=33.6e-15 PD=760e-9 PS=760e-9 NRD=1.16667 NRS=1.16667 M=1
mi0__i3__nm0 n12__i0__i3__net1 n2__i0__net1 n3__i0__net8 n3__vss g45n1svt L=45e-9 W=120e-9 AD=16.8e-15 AS=16.8e-15 PD=520e-9 PS=520e-9 NRD=1.16667 NRS=1.16667 M=1
mi0__i3__nm8 n127__vss n2__i0__i3__net2 n8__i0__i3__net1 n3__vss g45n1svt L=570e-9 W=120e-9 AD=16.8e-15 AS=16.8e-15 PD=520e-9 PS=520e-9 NRD=1.16667 NRS=1.16667 M=1
mi0__i3__nm18 n124__vss n7__rst n15__i0__i3__net1 n3__vss g45n1svt L=45e-9 W=120e-9 AD=16.8e-15 AS=16.8e-15 PD=520e-9 PS=520e-9 NRD=1.16667 NRS=1.16667 M=1
mi0__i3__nm2_1__rcx n9__i0__i3__net2 n6__i0__i3__net1 n122__vss n3__vss g45n1svt L=45e-9 W=240e-9 AD=38.4e-15 AS=38.4e-15 PD=780e-9 PS=780e-9 NRD=1.16667 NRS=1.16667 M=1
mi0__i3__nm2 n121__vss n5__i0__i3__net1 n9__i0__i3__net2 n3__vss g45n1svt L=45e-9 W=240e-9 AD=33.6e-15 AS=33.6e-15 PD=780e-9 PS=780e-9 NRD=1.16667 NRS=1.16667 M=1
mi0__i3__nm12 n12__i0__i3__net5 n4__i0__net7 n10__i0__i3__net2 n3__vss g45n1svt L=45e-9 W=120e-9 AD=16.8e-15 AS=16.8e-15 PD=520e-9 PS=520e-9 NRD=1.16667 NRS=1.16667 M=1
mi0__i3__nm15 n118__vss n2__i0__i3__net4 n8__i0__i3__net5 n3__vss g45n1svt L=570e-9 W=120e-9 AD=16.8e-15 AS=16.8e-15 PD=520e-9 PS=520e-9 NRD=1.16667 NRS=1.16667 M=1
mi0__i3__nm13_1__rcx n8__i0__i3__net4 n6__i0__i3__net5 n116__vss n3__vss g45n1svt L=45e-9 W=240e-9 AD=38.4e-15 AS=38.4e-15 PD=780e-9 PS=780e-9 NRD=1.16667 NRS=1.16667 M=1
mi0__i3__nm13 n114__vss n5__i0__i3__net5 n8__i0__i3__net4 n3__vss g45n1svt L=45e-9 W=240e-9 AD=33.6e-15 AS=33.6e-15 PD=780e-9 PS=780e-9 NRD=1.16667 NRS=1.16667 M=1
mi0__i3__nm16 n20__i0__net8 n6__i0__i3__net4 n113__vss n3__vss g45n1svt L=45e-9 W=240e-9 AD=33.6e-15 AS=33.6e-15 PD=760e-9 PS=760e-9 NRD=1.16667 NRS=1.16667 M=1
mi0__i3__nm17 n12__i0__net11 n9__i0__net8 n111__vss n3__vss g45n1svt L=45e-9 W=240e-9 AD=33.6e-15 AS=33.6e-15 PD=760e-9 PS=760e-9 NRD=1.16667 NRS=1.16667 M=1
mi0__i4__nm3 n10__i0__net9 n3__i0__net11 n108__vss n3__vss g45n1svt L=45e-9 W=120e-9 AD=19.2e-15 AS=19.2e-15 PD=540e-9 PS=540e-9 NRD=1.16667 NRS=1.16667 M=1
mi0__i4__nm2 n57__vdd n13__i0__net8 n10__i0__net9 n3__vss g45n1svt L=45e-9 W=120e-9 AD=16.8e-15 AS=16.8e-15 PD=540e-9 PS=540e-9 NRD=1.16667 NRS=1.16667 M=1
mi0__i4__nm6 n11__i0__net10 n7__i0__net9 n107__vss n3__vss g45n1svt L=45e-9 W=240e-9 AD=33.6e-15 AS=33.6e-15 PD=760e-9 PS=760e-9 NRD=1.16667 NRS=1.16667 M=1
mi0__i4__nm5 n104__vss n7__i0__net10 n18__i0__net9 n3__vss g45n1svt L=45e-9 W=240e-9 AD=33.6e-15 AS=33.6e-15 PD=760e-9 PS=760e-9 NRD=1.16667 NRS=1.16667 M=1
mi0__i4__nm1 n18__i0__net10 n4__i0__net11 n43__vdd n3__vss g45n1svt L=45e-9 W=120e-9 AD=19.2e-15 AS=19.2e-15 PD=540e-9 PS=540e-9 NRD=1.16667 NRS=1.16667 M=1
mi0__i4__nm0 n100__vss n14__i0__net8 n18__i0__net10 n3__vss g45n1svt L=45e-9 W=120e-9 AD=16.8e-15 AS=16.8e-15 PD=540e-9 PS=540e-9 NRD=1.16667 NRS=1.16667 M=1
mi0__nm0 n5__i0__net3 n1__clk n46__vss n3__vss g45n1svt L=45e-9 W=120e-9 AD=16.8e-15 AS=16.8e-15 PD=520e-9 PS=520e-9 NRD=1.16667 NRS=1.16667 M=1
mi0__nm1 n7__i0__net6 n3__rst n129__vss n3__vss g45n1svt L=45e-9 W=120e-9 AD=16.8e-15 AS=16.8e-15 PD=520e-9 PS=520e-9 NRD=1.16667 NRS=1.16667 M=1
mi0__nm14 n25__net11 i0__net10 n24__vss n3__vss g45n1svt L=45e-9 W=240e-9 AD=33.6e-15 AS=33.6e-15 PD=760e-9 PS=760e-9 NRD=1.16667 NRS=1.16667 M=1
mi0__nm15 n26__net7 i0__net9 n22__vss n3__vss g45n1svt L=45e-9 W=240e-9 AD=33.6e-15 AS=33.6e-15 PD=760e-9 PS=760e-9 NRD=1.16667 NRS=1.16667 M=1
mi7__nm0 n13__i7__net1 n34__net9 n3__y_in_3 n3__vss g45n1svt L=45e-9 W=120e-9 AD=16.8e-15 AS=16.8e-15 PD=520e-9 PS=520e-9 NRD=1.16667 NRS=1.16667 M=1
mi7__nm8 n106__vss n3__i7__net2 n8__i7__net1 n3__vss g45n1svt L=570e-9 W=120e-9 AD=16.8e-15 AS=16.8e-15 PD=520e-9 PS=520e-9 NRD=1.16667 NRS=1.16667 M=1
mi7__nm18 n105__vss n30__net3 n15__i7__net1 n3__vss g45n1svt L=45e-9 W=120e-9 AD=16.8e-15 AS=16.8e-15 PD=520e-9 PS=520e-9 NRD=1.16667 NRS=1.16667 M=1
mi7__nm2_1__rcx n11__i7__net2 n7__i7__net1 n103__vss n3__vss g45n1svt L=45e-9 W=240e-9 AD=38.4e-15 AS=38.4e-15 PD=780e-9 PS=780e-9 NRD=1.16667 NRS=1.16667 M=1
mi7__nm2 n102__vss i7__net1 n11__i7__net2 n3__vss g45n1svt L=45e-9 W=240e-9 AD=33.6e-15 AS=33.6e-15 PD=780e-9 PS=780e-9 NRD=1.16667 NRS=1.16667 M=1
mi7__nm12 n13__i7__net5 n58__net10 n5__i7__net2 n3__vss g45n1svt L=45e-9 W=120e-9 AD=16.8e-15 AS=16.8e-15 PD=520e-9 PS=520e-9 NRD=1.16667 NRS=1.16667 M=1
mi7__nm15 n96__vss n3__i7__net4 n8__i7__net5 n3__vss g45n1svt L=570e-9 W=120e-9 AD=16.8e-15 AS=16.8e-15 PD=520e-9 PS=520e-9 NRD=1.16667 NRS=1.16667 M=1
mi7__nm13_1__rcx n8__i7__net4 n7__i7__net5 n94__vss n3__vss g45n1svt L=45e-9 W=240e-9 AD=38.4e-15 AS=38.4e-15 PD=780e-9 PS=780e-9 NRD=1.16667 NRS=1.16667 M=1
mi7__nm13 n92__vss i7__net5 n8__i7__net4 n3__vss g45n1svt L=45e-9 W=240e-9 AD=33.6e-15 AS=33.6e-15 PD=780e-9 PS=780e-9 NRD=1.16667 NRS=1.16667 M=1
mi7__nm16 n8__y_out_b_3 n4__i7__net4 n90__vss n3__vss g45n1svt L=45e-9 W=240e-9 AD=33.6e-15 AS=33.6e-15 PD=760e-9 PS=760e-9 NRD=1.16667 NRS=1.16667 M=1
mi7__nm17 n1__y_out_3 n1__y_out_b_3 n88__vss n3__vss g45n1svt L=45e-9 W=240e-9 AD=33.6e-15 AS=33.6e-15 PD=760e-9 PS=760e-9 NRD=1.16667 NRS=1.16667 M=1
mi1__nm0 n13__i1__net1 n2__net9 n1__x_in_3 n3__vss g45n1svt L=45e-9 W=120e-9 AD=16.8e-15 AS=16.8e-15 PD=520e-9 PS=520e-9 NRD=1.16667 NRS=1.16667 M=1
mi1__nm8 n128__vss n3__i1__net2 n8__i1__net1 n3__vss g45n1svt L=570e-9 W=120e-9 AD=16.8e-15 AS=16.8e-15 PD=520e-9 PS=520e-9 NRD=1.16667 NRS=1.16667 M=1
mi1__nm18 n126__vss n2__net3 n15__i1__net1 n3__vss g45n1svt L=45e-9 W=120e-9 AD=16.8e-15 AS=16.8e-15 PD=520e-9 PS=520e-9 NRD=1.16667 NRS=1.16667 M=1
mi1__nm2_1__rcx n12__i1__net2 n7__i1__net1 n125__vss n3__vss g45n1svt L=45e-9 W=240e-9 AD=38.4e-15 AS=38.4e-15 PD=780e-9 PS=780e-9 NRD=1.16667 NRS=1.16667 M=1
mi1__nm2 n123__vss i1__net1 n12__i1__net2 n3__vss g45n1svt L=45e-9 W=240e-9 AD=33.6e-15 AS=33.6e-15 PD=780e-9 PS=780e-9 NRD=1.16667 NRS=1.16667 M=1
mi1__nm12 n13__i1__net5 n10__net10 n6__i1__net2 n3__vss g45n1svt L=45e-9 W=120e-9 AD=16.8e-15 AS=16.8e-15 PD=520e-9 PS=520e-9 NRD=1.16667 NRS=1.16667 M=1
mi1__nm15 n120__vss n3__i1__net4 n8__i1__net5 n3__vss g45n1svt L=570e-9 W=120e-9 AD=16.8e-15 AS=16.8e-15 PD=520e-9 PS=520e-9 NRD=1.16667 NRS=1.16667 M=1
mi1__nm13_1__rcx n8__i1__net4 n7__i1__net5 n119__vss n3__vss g45n1svt L=45e-9 W=240e-9 AD=38.4e-15 AS=38.4e-15 PD=780e-9 PS=780e-9 NRD=1.16667 NRS=1.16667 M=1
mi1__nm13 n117__vss i1__net5 n8__i1__net4 n3__vss g45n1svt L=45e-9 W=240e-9 AD=33.6e-15 AS=33.6e-15 PD=780e-9 PS=780e-9 NRD=1.16667 NRS=1.16667 M=1
mi1__nm16 n8__x_out_b_3 n4__i1__net4 n115__vss n3__vss g45n1svt L=45e-9 W=240e-9 AD=33.6e-15 AS=33.6e-15 PD=760e-9 PS=760e-9 NRD=1.16667 NRS=1.16667 M=1
mi1__nm17 n1__x_out_3 n1__x_out_b_3 n112__vss n3__vss g45n1svt L=45e-9 W=240e-9 AD=33.6e-15 AS=33.6e-15 PD=760e-9 PS=760e-9 NRD=1.16667 NRS=1.16667 M=1
mi4__nm0 n13__i4__net1 n38__net9 n3__y_in_1 n3__vss g45n1svt L=45e-9 W=120e-9 AD=16.8e-15 AS=16.8e-15 PD=520e-9 PS=520e-9 NRD=1.16667 NRS=1.16667 M=1
mi4__nm8 n170__vss n3__i4__net2 n8__i4__net1 n3__vss g45n1svt L=570e-9 W=120e-9 AD=16.8e-15 AS=16.8e-15 PD=520e-9 PS=520e-9 NRD=1.16667 NRS=1.16667 M=1
mi4__nm18 n168__vss n34__net3 n15__i4__net1 n3__vss g45n1svt L=45e-9 W=120e-9 AD=16.8e-15 AS=16.8e-15 PD=520e-9 PS=520e-9 NRD=1.16667 NRS=1.16667 M=1
mi4__nm2_1__rcx n11__i4__net2 n7__i4__net1 n166__vss n3__vss g45n1svt L=45e-9 W=240e-9 AD=38.4e-15 AS=38.4e-15 PD=780e-9 PS=780e-9 NRD=1.16667 NRS=1.16667 M=1
mi4__nm2 n164__vss i4__net1 n11__i4__net2 n3__vss g45n1svt L=45e-9 W=240e-9 AD=33.6e-15 AS=33.6e-15 PD=780e-9 PS=780e-9 NRD=1.16667 NRS=1.16667 M=1
mi4__nm12 n13__i4__net5 n62__net10 n5__i4__net2 n3__vss g45n1svt L=45e-9 W=120e-9 AD=16.8e-15 AS=16.8e-15 PD=520e-9 PS=520e-9 NRD=1.16667 NRS=1.16667 M=1
mi4__nm15 n162__vss n3__i4__net4 n8__i4__net5 n3__vss g45n1svt L=570e-9 W=120e-9 AD=16.8e-15 AS=16.8e-15 PD=520e-9 PS=520e-9 NRD=1.16667 NRS=1.16667 M=1
mi4__nm13_1__rcx n8__i4__net4 n7__i4__net5 n160__vss n3__vss g45n1svt L=45e-9 W=240e-9 AD=38.4e-15 AS=38.4e-15 PD=780e-9 PS=780e-9 NRD=1.16667 NRS=1.16667 M=1
mi4__nm13 n158__vss i4__net5 n8__i4__net4 n3__vss g45n1svt L=45e-9 W=240e-9 AD=33.6e-15 AS=33.6e-15 PD=780e-9 PS=780e-9 NRD=1.16667 NRS=1.16667 M=1
mi4__nm16 n8__y_out_b_1 n4__i4__net4 n156__vss n3__vss g45n1svt L=45e-9 W=240e-9 AD=33.6e-15 AS=33.6e-15 PD=760e-9 PS=760e-9 NRD=1.16667 NRS=1.16667 M=1
mi4__nm17 n1__y_out_1 n1__y_out_b_1 n155__vss n3__vss g45n1svt L=45e-9 W=240e-9 AD=33.6e-15 AS=33.6e-15 PD=760e-9 PS=760e-9 NRD=1.16667 NRS=1.16667 M=1
mi3__nm0 n13__i3__net1 n6__net9 n1__x_in_1 n3__vss g45n1svt L=45e-9 W=120e-9 AD=16.8e-15 AS=16.8e-15 PD=520e-9 PS=520e-9 NRD=1.16667 NRS=1.16667 M=1
mi3__nm8 n188__vss n3__i3__net2 n8__i3__net1 n3__vss g45n1svt L=570e-9 W=120e-9 AD=16.8e-15 AS=16.8e-15 PD=520e-9 PS=520e-9 NRD=1.16667 NRS=1.16667 M=1
mi3__nm18 n186__vss n6__net3 n15__i3__net1 n3__vss g45n1svt L=45e-9 W=120e-9 AD=16.8e-15 AS=16.8e-15 PD=520e-9 PS=520e-9 NRD=1.16667 NRS=1.16667 M=1
mi3__nm2_1__rcx n12__i3__net2 n7__i3__net1 n184__vss n3__vss g45n1svt L=45e-9 W=240e-9 AD=38.4e-15 AS=38.4e-15 PD=780e-9 PS=780e-9 NRD=1.16667 NRS=1.16667 M=1
mi3__nm2 n182__vss i3__net1 n12__i3__net2 n3__vss g45n1svt L=45e-9 W=240e-9 AD=33.6e-15 AS=33.6e-15 PD=780e-9 PS=780e-9 NRD=1.16667 NRS=1.16667 M=1
mi3__nm12 n13__i3__net5 n14__net10 n6__i3__net2 n3__vss g45n1svt L=45e-9 W=120e-9 AD=16.8e-15 AS=16.8e-15 PD=520e-9 PS=520e-9 NRD=1.16667 NRS=1.16667 M=1
mi3__nm15 n180__vss n3__i3__net4 n8__i3__net5 n3__vss g45n1svt L=570e-9 W=120e-9 AD=16.8e-15 AS=16.8e-15 PD=520e-9 PS=520e-9 NRD=1.16667 NRS=1.16667 M=1
mi3__nm13_1__rcx n8__i3__net4 n7__i3__net5 n178__vss n3__vss g45n1svt L=45e-9 W=240e-9 AD=38.4e-15 AS=38.4e-15 PD=780e-9 PS=780e-9 NRD=1.16667 NRS=1.16667 M=1
mi3__nm13 n176__vss i3__net5 n8__i3__net4 n3__vss g45n1svt L=45e-9 W=240e-9 AD=33.6e-15 AS=33.6e-15 PD=780e-9 PS=780e-9 NRD=1.16667 NRS=1.16667 M=1
mi3__nm16 n8__x_out_b_1 n4__i3__net4 n174__vss n3__vss g45n1svt L=45e-9 W=240e-9 AD=33.6e-15 AS=33.6e-15 PD=760e-9 PS=760e-9 NRD=1.16667 NRS=1.16667 M=1
mi3__nm17 n1__x_out_1 n1__x_out_b_1 n172__vss n3__vss g45n1svt L=45e-9 W=240e-9 AD=33.6e-15 AS=33.6e-15 PD=760e-9 PS=760e-9 NRD=1.16667 NRS=1.16667 M=1
mi6__nm0 n12__i6__net1 n36__net9 n5__y_in_2 n3__vss g45n1svt L=45e-9 W=120e-9 AD=16.8e-15 AS=16.8e-15 PD=520e-9 PS=520e-9 NRD=1.16667 NRS=1.16667 M=1
mi6__nm8 n171__vss n2__i6__net2 n8__i6__net1 n3__vss g45n1svt L=570e-9 W=120e-9 AD=16.8e-15 AS=16.8e-15 PD=520e-9 PS=520e-9 NRD=1.16667 NRS=1.16667 M=1
mi6__nm18 n169__vss n32__net3 n15__i6__net1 n3__vss g45n1svt L=45e-9 W=120e-9 AD=16.8e-15 AS=16.8e-15 PD=520e-9 PS=520e-9 NRD=1.16667 NRS=1.16667 M=1
mi6__nm2_1__rcx n8__i6__net2 n6__i6__net1 n167__vss n3__vss g45n1svt L=45e-9 W=240e-9 AD=38.4e-15 AS=38.4e-15 PD=780e-9 PS=780e-9 NRD=1.16667 NRS=1.16667 M=1
mi6__nm2 n165__vss n5__i6__net1 n8__i6__net2 n3__vss g45n1svt L=45e-9 W=240e-9 AD=33.6e-15 AS=33.6e-15 PD=780e-9 PS=780e-9 NRD=1.16667 NRS=1.16667 M=1
mi6__nm12 n12__i6__net5 n60__net10 n9__i6__net2 n3__vss g45n1svt L=45e-9 W=120e-9 AD=16.8e-15 AS=16.8e-15 PD=520e-9 PS=520e-9 NRD=1.16667 NRS=1.16667 M=1
mi6__nm15 n163__vss n2__i6__net4 n8__i6__net5 n3__vss g45n1svt L=570e-9 W=120e-9 AD=16.8e-15 AS=16.8e-15 PD=520e-9 PS=520e-9 NRD=1.16667 NRS=1.16667 M=1
mi6__nm13_1__rcx n8__i6__net4 n6__i6__net5 n161__vss n3__vss g45n1svt L=45e-9 W=240e-9 AD=38.4e-15 AS=38.4e-15 PD=780e-9 PS=780e-9 NRD=1.16667 NRS=1.16667 M=1
mi6__nm13 n159__vss n5__i6__net5 n8__i6__net4 n3__vss g45n1svt L=45e-9 W=240e-9 AD=33.6e-15 AS=33.6e-15 PD=780e-9 PS=780e-9 NRD=1.16667 NRS=1.16667 M=1
mi6__nm16 n6__y_out_b_2 n6__i6__net4 n157__vss n3__vss g45n1svt L=45e-9 W=240e-9 AD=33.6e-15 AS=33.6e-15 PD=760e-9 PS=760e-9 NRD=1.16667 NRS=1.16667 M=1
mi6__nm17 n3__y_out_2 n4__y_out_b_2 n131__vss n3__vss g45n1svt L=45e-9 W=240e-9 AD=33.6e-15 AS=33.6e-15 PD=760e-9 PS=760e-9 NRD=1.16667 NRS=1.16667 M=1
mi2__nm0 n12__i2__net1 n4__net9 n3__x_in_2 n3__vss g45n1svt L=45e-9 W=120e-9 AD=16.8e-15 AS=16.8e-15 PD=520e-9 PS=520e-9 NRD=1.16667 NRS=1.16667 M=1
mi2__nm8 n189__vss n2__i2__net2 n8__i2__net1 n3__vss g45n1svt L=570e-9 W=120e-9 AD=16.8e-15 AS=16.8e-15 PD=520e-9 PS=520e-9 NRD=1.16667 NRS=1.16667 M=1
mi2__nm18 n187__vss n4__net3 n15__i2__net1 n3__vss g45n1svt L=45e-9 W=120e-9 AD=16.8e-15 AS=16.8e-15 PD=520e-9 PS=520e-9 NRD=1.16667 NRS=1.16667 M=1
mi2__nm2_1__rcx n9__i2__net2 n6__i2__net1 n185__vss n3__vss g45n1svt L=45e-9 W=240e-9 AD=38.4e-15 AS=38.4e-15 PD=780e-9 PS=780e-9 NRD=1.16667 NRS=1.16667 M=1
mi2__nm2 n183__vss n5__i2__net1 n9__i2__net2 n3__vss g45n1svt L=45e-9 W=240e-9 AD=33.6e-15 AS=33.6e-15 PD=780e-9 PS=780e-9 NRD=1.16667 NRS=1.16667 M=1
mi2__nm12 n12__i2__net5 n12__net10 n10__i2__net2 n3__vss g45n1svt L=45e-9 W=120e-9 AD=16.8e-15 AS=16.8e-15 PD=520e-9 PS=520e-9 NRD=1.16667 NRS=1.16667 M=1
mi2__nm15 n181__vss n2__i2__net4 n8__i2__net5 n3__vss g45n1svt L=570e-9 W=120e-9 AD=16.8e-15 AS=16.8e-15 PD=520e-9 PS=520e-9 NRD=1.16667 NRS=1.16667 M=1
mi2__nm13_1__rcx n8__i2__net4 n6__i2__net5 n179__vss n3__vss g45n1svt L=45e-9 W=240e-9 AD=38.4e-15 AS=38.4e-15 PD=780e-9 PS=780e-9 NRD=1.16667 NRS=1.16667 M=1
mi2__nm13 n177__vss n5__i2__net5 n8__i2__net4 n3__vss g45n1svt L=45e-9 W=240e-9 AD=33.6e-15 AS=33.6e-15 PD=780e-9 PS=780e-9 NRD=1.16667 NRS=1.16667 M=1
mi2__nm16 n6__x_out_b_2 n6__i2__net4 n175__vss n3__vss g45n1svt L=45e-9 W=240e-9 AD=33.6e-15 AS=33.6e-15 PD=760e-9 PS=760e-9 NRD=1.16667 NRS=1.16667 M=1
mi2__nm17 n3__x_out_2 n4__x_out_b_2 n173__vss n3__vss g45n1svt L=45e-9 W=240e-9 AD=33.6e-15 AS=33.6e-15 PD=760e-9 PS=760e-9 NRD=1.16667 NRS=1.16667 M=1
mi5__nm0 n12__i5__net1 n40__net9 n5__y_in_0 n3__vss g45n1svt L=45e-9 W=120e-9 AD=16.8e-15 AS=16.8e-15 PD=520e-9 PS=520e-9 NRD=1.16667 NRS=1.16667 M=1
mi5__nm8 n220__vss n2__i5__net2 n8__i5__net1 n3__vss g45n1svt L=570e-9 W=120e-9 AD=16.8e-15 AS=16.8e-15 PD=520e-9 PS=520e-9 NRD=1.16667 NRS=1.16667 M=1
mi5__nm18 n219__vss n36__net3 n15__i5__net1 n3__vss g45n1svt L=45e-9 W=120e-9 AD=16.8e-15 AS=16.8e-15 PD=520e-9 PS=520e-9 NRD=1.16667 NRS=1.16667 M=1
mi5__nm2_1__rcx n8__i5__net2 n6__i5__net1 n218__vss n3__vss g45n1svt L=45e-9 W=240e-9 AD=38.4e-15 AS=38.4e-15 PD=780e-9 PS=780e-9 NRD=1.16667 NRS=1.16667 M=1
mi5__nm2 n217__vss n5__i5__net1 n8__i5__net2 n3__vss g45n1svt L=45e-9 W=240e-9 AD=33.6e-15 AS=33.6e-15 PD=780e-9 PS=780e-9 NRD=1.16667 NRS=1.16667 M=1
mi5__nm12 n12__i5__net5 n64__net10 n9__i5__net2 n3__vss g45n1svt L=45e-9 W=120e-9 AD=16.8e-15 AS=16.8e-15 PD=520e-9 PS=520e-9 NRD=1.16667 NRS=1.16667 M=1
mi5__nm15 n216__vss n2__i5__net4 n8__i5__net5 n3__vss g45n1svt L=570e-9 W=120e-9 AD=16.8e-15 AS=16.8e-15 PD=520e-9 PS=520e-9 NRD=1.16667 NRS=1.16667 M=1
mi5__nm13_1__rcx n8__i5__net4 n6__i5__net5 n215__vss n3__vss g45n1svt L=45e-9 W=240e-9 AD=38.4e-15 AS=38.4e-15 PD=780e-9 PS=780e-9 NRD=1.16667 NRS=1.16667 M=1
mi5__nm13 n214__vss n5__i5__net5 n8__i5__net4 n3__vss g45n1svt L=45e-9 W=240e-9 AD=33.6e-15 AS=33.6e-15 PD=780e-9 PS=780e-9 NRD=1.16667 NRS=1.16667 M=1
mi5__nm16 n6__y_out_b_0 n6__i5__net4 n213__vss n3__vss g45n1svt L=45e-9 W=240e-9 AD=33.6e-15 AS=33.6e-15 PD=760e-9 PS=760e-9 NRD=1.16667 NRS=1.16667 M=1
mi5__nm17 n3__y_out_0 n4__y_out_b_0 n190__vss n3__vss g45n1svt L=45e-9 W=240e-9 AD=33.6e-15 AS=33.6e-15 PD=760e-9 PS=760e-9 NRD=1.16667 NRS=1.16667 M=1
mi8__nm0 n12__i8__net1 n8__net9 n3__x_in_0 n3__vss g45n1svt L=45e-9 W=120e-9 AD=16.8e-15 AS=16.8e-15 PD=520e-9 PS=520e-9 NRD=1.16667 NRS=1.16667 M=1
mi8__nm8 n229__vss n2__i8__net2 n8__i8__net1 n3__vss g45n1svt L=570e-9 W=120e-9 AD=16.8e-15 AS=16.8e-15 PD=520e-9 PS=520e-9 NRD=1.16667 NRS=1.16667 M=1
mi8__nm18 n228__vss n8__net3 n15__i8__net1 n3__vss g45n1svt L=45e-9 W=120e-9 AD=16.8e-15 AS=16.8e-15 PD=520e-9 PS=520e-9 NRD=1.16667 NRS=1.16667 M=1
mi8__nm2_1__rcx n9__i8__net2 n6__i8__net1 n227__vss n3__vss g45n1svt L=45e-9 W=240e-9 AD=38.4e-15 AS=38.4e-15 PD=780e-9 PS=780e-9 NRD=1.16667 NRS=1.16667 M=1
mi8__nm2 n226__vss n5__i8__net1 n9__i8__net2 n3__vss g45n1svt L=45e-9 W=240e-9 AD=33.6e-15 AS=33.6e-15 PD=780e-9 PS=780e-9 NRD=1.16667 NRS=1.16667 M=1
mi8__nm12 n12__i8__net5 n16__net10 n10__i8__net2 n3__vss g45n1svt L=45e-9 W=120e-9 AD=16.8e-15 AS=16.8e-15 PD=520e-9 PS=520e-9 NRD=1.16667 NRS=1.16667 M=1
mi8__nm15 n225__vss n2__i8__net4 n8__i8__net5 n3__vss g45n1svt L=570e-9 W=120e-9 AD=16.8e-15 AS=16.8e-15 PD=520e-9 PS=520e-9 NRD=1.16667 NRS=1.16667 M=1
mi8__nm13_1__rcx n8__i8__net4 n6__i8__net5 n224__vss n3__vss g45n1svt L=45e-9 W=240e-9 AD=38.4e-15 AS=38.4e-15 PD=780e-9 PS=780e-9 NRD=1.16667 NRS=1.16667 M=1
mi8__nm13 n223__vss n5__i8__net5 n8__i8__net4 n3__vss g45n1svt L=45e-9 W=240e-9 AD=33.6e-15 AS=33.6e-15 PD=780e-9 PS=780e-9 NRD=1.16667 NRS=1.16667 M=1
mi8__nm16 n6__x_out_b_0 n6__i8__net4 n222__vss n3__vss g45n1svt L=45e-9 W=240e-9 AD=33.6e-15 AS=33.6e-15 PD=760e-9 PS=760e-9 NRD=1.16667 NRS=1.16667 M=1
mi8__nm17 n3__x_out_0 n4__x_out_b_0 n221__vss n3__vss g45n1svt L=45e-9 W=240e-9 AD=33.6e-15 AS=33.6e-15 PD=760e-9 PS=760e-9 NRD=1.16667 NRS=1.16667 M=1
mnm10 n2__clk_div4_out_b net7 n13__vss n3__vss g45n1svt L=45e-9 W=240e-9 AD=33.6e-15 AS=33.6e-15 PD=760e-9 PS=760e-9 NRD=1.16667 NRS=1.16667 M=1
mnm9 n1__clk_div4_out net11 n12__vss n3__vss g45n1svt L=45e-9 W=240e-9 AD=33.6e-15 AS=33.6e-15 PD=760e-9 PS=760e-9 NRD=1.16667 NRS=1.16667 M=1


cxo0  x_out_0   vss 2f
cxo1  x_out_1   vss 2f
cxo2  x_out_2   vss 2f
cxo3  x_out_3   vss 2f
cxob0 x_out_b_0 vss 2f
cxob1 x_out_b_1 vss 2f
cxob2 x_out_b_2 vss 2f
cxob3 x_out_b_3 vss 2f
cyo0  y_out_0   vss 2f
cyo1  y_out_1   vss 2f
cyo2  y_out_2   vss 2f
cyo3  y_out_3   vss 2f
cyob0 y_out_b_0 vss 2f
cyob1 y_out_b_1 vss 2f
cyob2 y_out_b_2 vss 2f
cyob3 y_out_b_3 vss 2f

cclk_out   clk_div4_out   vss 0.66f
cclk_out_b clk_div4_out_b vss 0.66f

.ends data_reg_bank