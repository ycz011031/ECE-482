.subckt Top_Level CK Reset x0 x1 x2 x3 y0 y1 y2 y3 Serial_out R_OUT vddio vdd vss

c1 vdd vss 3.361e-15
c2 ck vss 168.261e-18
c3 reset vss 203.737e-18
c4 x0 vss 9.60712e-18
c5 x1 vss 8.96121e-18
c6 x2 vss 9.60712e-18
c7 x3 vss 8.98678e-18
c8 y0 vss 227.549e-18
c9 y1 vss 279.82e-18
c10 y2 vss 279.832e-18
c11 y3 vss 242.187e-18
c12 r_out vss 1.06173e-15
c13 serial_out vss 49.6725e-18
c14 vddio vss 1.58567e-15
c15 serial_out_b_high vss 53.116e-18
c16 serial_out_b_high_buff vss 75.0592e-18
c17 ck4 vss 93.2156e-18
c18 reset_b vss 17.7248e-18
c19 shift vss 33.3982e-18
c20 reset_buff vss 21.8848e-18
c21 ck_b vss 28.9096e-18
c22 ck_buff vss 26.5674e-18
c23 y_out_2 vss 18.5219e-18
c24 x_out_1 vss 56.1667e-18
c25 y_out_1 vss 23.679e-18
c26 x_out_3 vss 50.386e-18
c27 y_out_3 vss 21.2741e-18
c28 r0 vss 104.731e-18
c29 r1 vss 26.3309e-18
c30 r2 vss 36.4124e-18
c31 y_out_0 vss 19.4176e-18
c32 x_out_0 vss 97.3253e-18
c33 x_out_2 vss 97.3253e-18
c34 r2_buff vss 171.829e-18
c35 net3 vss 71.8655e-18
c36 r1_buff vss 240.131e-18
c37 net4 vss 53.836e-18
c38 r0_buff vss 196.842e-18
c39 net8 vss 21.6782e-18
c40 net7 vss 19.2528e-18
c41 net14 vss 21.8468e-18
c42 net10 vss 50.0994e-18
c43 net6 vss 20.3954e-18
c44 net9 vss 68.8515e-18
c45 net13 vss 13.8799e-18
c46 i2__q vss 69.2281e-18
c47 i2__net76 vss 21.1694e-18
c48 i2__net73 vss 75.7598e-18
c49 i2__net1 vss 31.6483e-18
c50 i2__net77 vss 114.292e-18
c51 i2__net74 vss 24.8938e-18
c52 i2__net75 vss 113.256e-18
c53 i2__net79 vss 31.8761e-18
c54 i1__q vss 46.539e-18
c55 i1__net76 vss 18.6724e-18
c56 i1__net73 vss 25.3983e-18
c57 i1__net1 vss 22.7684e-18
c58 i1__net77 vss 117.54e-18
c59 i1__net74 vss 19.1442e-18
c60 i1__net75 vss 119.711e-18
c61 i1__net79 vss 31.1634e-18
c62 i0__q vss 76.4322e-18
c63 i0__net76 vss 24.0399e-18
c64 i0__net73 vss 80.3364e-18
c65 i0__net1 vss 30.2825e-18
c66 i0__net77 vss 112.046e-18
c67 i0__net74 vss 26.531e-18
c68 i0__net75 vss 112.56e-18
c69 i0__net79 vss 32.0412e-18
c70 i14__clk_div4_out_b vss 156.249e-18
c71 i14__net7 vss 20.305e-18
c72 i14__net11 vss 22.3205e-18
c73 i14__net9 vss 31.6438e-18
c74 i14__x_out_b_3 vss 30.4937e-18
c75 i14__net10 vss 29.561e-18
c76 i14__net3 vss 21.4174e-18
c77 i14__net4 vss 16.5107e-18
c78 i14__x_out_b_0 vss 28.9656e-18
c79 i14__y_out_b_0 vss 30.4937e-18
c80 i14__y_out_b_2 vss 28.0669e-18
c81 i14__x_out_b_2 vss 21.8154e-18
c82 i14__y_out_b_1 vss 22.7404e-18
c83 i14__y_out_b_3 vss 24.1155e-18
c84 i14__x_out_b_1 vss 21.3989e-18
c85 i3__avs50 vss 197.088e-18
c86 i14__i17__net10 vss 21.6249e-18
c87 i14__i17__net9 vss 22.1197e-18
c88 i14__i17__net8 vss 58.4991e-18
c89 i14__i17__net11 vss 32.7911e-18
c90 i14__i17__net1 vss 31.1122e-18
c91 i14__i17__net7 vss 28.5496e-18
c92 i14__i17__net6 vss 16.3976e-18
c93 i14__i17__net3 vss 28.9417e-18
c94 i14__i17__i2__net5 vss 17.4278e-18
c95 i14__i17__i2__net4 vss 116.515e-18
c96 i14__i17__i2__net1 vss 17.1811e-18
c97 i14__i17__i2__net2 vss 116.758e-18
c98 i14__i17__i3__net5 vss 24.8353e-18
c99 i14__i17__i3__net4 vss 112.457e-18
c100 i14__i17__i3__net1 vss 26.5256e-18
c101 i14__i17__i3__net2 vss 113.265e-18
c102 i14__i11__net5 vss 19.924e-18
c103 i14__i11__net4 vss 119.199e-18
c104 i14__i11__net1 vss 21.8584e-18
c105 i14__i11__net2 vss 118.31e-18
c106 i14__i13__net5 vss 18.9608e-18
c107 i14__i13__net4 vss 116.762e-18
c108 i14__i13__net1 vss 20.2696e-18
c109 i14__i13__net2 vss 118.427e-18
c110 i14__i15__net5 vss 18.5487e-18
c111 i14__i15__net4 vss 116.339e-18
c112 i14__i15__net1 vss 18.8969e-18
c113 i14__i15__net2 vss 117.905e-18
c114 i14__i10__net5 vss 18.7278e-18
c115 i14__i10__net4 vss 115.551e-18
c116 i14__i10__net1 vss 19.4125e-18
c117 i14__i10__net2 vss 118.751e-18
c118 i14__i14__net5 vss 24.425e-18
c119 i14__i14__net4 vss 111.992e-18
c120 i14__i14__net1 vss 26.2874e-18
c121 i14__i14__net2 vss 111.764e-18
c122 i14__i16__net5 vss 24.0926e-18
c123 i14__i16__net4 vss 111.026e-18
c124 i14__i16__net1 vss 26.1676e-18
c125 i14__i16__net2 vss 112.527e-18
c126 i14__i12__net5 vss 24.4762e-18
c127 i14__i12__net4 vss 110.168e-18
c128 i14__i12__net1 vss 26.2901e-18
c129 i14__i12__net2 vss 111.258e-18
c130 i14__i9__net5 vss 24.0926e-18
c131 i14__i9__net4 vss 110.526e-18
c132 i14__i9__net1 vss 26.1676e-18
c133 i14__i9__net2 vss 112.42e-18
c134 i13__net3 vss 25.651e-18
c135 i13__net23 vss 48.6792e-18
c136 i13__net17 vss 39.5137e-18
c137 i13__a0 vss 44.5296e-18
c138 i13__a1 vss 33.549e-18
c139 i13__a2 vss 31.5223e-18
c140 i13__a3 vss 41.1745e-18
c141 i13__net1 vss 35.1513e-18
c142 i13__net2 vss 43.6249e-18
c143 i13__net12 vss 34.1859e-18
c144 i13__net7 vss 45.5625e-18
c145 i13__net11 vss 40.9503e-18
c146 i13__net18 vss 32.5957e-18
c147 i13__i20__net3 vss 85.9308e-18
c148 i13__i20__net1 vss 26.4676e-18
c149 i13__i20__i4__net2 vss 18.0023e-18
c150 i13__i19__net3 vss 87.7249e-18
c151 i13__i19__net1 vss 23.8145e-18
c152 i13__i19__i4__net2 vss 20.6869e-18
c153 i13__i17__net3 vss 85.0196e-18
c154 i13__i17__net1 vss 25.0535e-18
c155 i13__i17__i4__net2 vss 19.7043e-18
c156 i13__i18__net3 vss 87.5787e-18
c157 i13__i18__net1 vss 26.6484e-18
c158 i13__i18__i4__net2 vss 20.5656e-18
c159 i13__i16__net3 vss 86.804e-18
c160 i13__i16__net1 vss 27.5924e-18
c161 i13__i16__i4__net2 vss 19.9575e-18
c162 i13__i15__net2 vss 19.1659e-18
c163 i13__i14__net2 vss 19.0016e-18
c164 i13__i13__net2 vss 20.4727e-18
c165 i13__i12__net2 vss 20.6068e-18
c166 i13__net6 vss 105.273e-18
c167 i9__net1 vss 28.5157e-18
c168 i9__i1__net1 vss 50.8258e-18
c169 i9__net2 vss 26.9181e-18
c170 i9__i4__net5 vss 22.1876e-18
c171 i9__i4__net4 vss 110.982e-18
c172 i9__i4__net1 vss 32.2288e-18
c173 i9__i4__net2 vss 110.506e-18
c174 i18__net5 vss 238.626e-18
c175 i18__net2 vss 144.241e-18
c176 i18__net1 vss 97.052e-18
c177 i18__net4 vss 229.458e-18
c178 i18__net3 vss 211.834e-18
c179 i12__bio vss 65.2048e-18
c180 i12__bcore_bar vss 139.122e-18
c181 n3__serial_out_b_high_buff vss 100.571e-18
c182 n5__serial_out_b_high vss 58.9234e-18
c183 n5__i18__net1 vss 109.027e-18
c184 n4__i18__net1 vss 117.27e-18
c185 n2__serial_out_b_high vss 53.5962e-18
c186 n7__i18__net2 vss 183.383e-18
c187 n8__i18__net2 vss 150.515e-18
c188 n10__i18__net2 vss 150.355e-18
c189 n2__i12__bio vss 47.5223e-18
c190 n6__i18__net2 vss 192.088e-18
c191 n30__i18__net3 vss 255.147e-18
c192 n27__i18__net3 vss 211.538e-18
c193 n24__i18__net3 vss 213.284e-18
c194 n21__i18__net3 vss 213.677e-18
c195 n18__i18__net3 vss 213.73e-18
c196 n15__i18__net3 vss 213.548e-18
c197 n12__i18__net3 vss 213.728e-18
c198 n9__i18__net3 vss 213.5e-18
c199 n6__i18__net3 vss 219.513e-18
c200 n3__i18__net3 vss 277.727e-18
c201 n122__i18__net4 vss 328.533e-18
c202 n115__i18__net4 vss 265.724e-18
c203 n112__i18__net4 vss 258.639e-18
c204 n105__i18__net4 vss 259.179e-18
c205 n102__i18__net4 vss 260.145e-18
c206 n97__i18__net4 vss 259.745e-18
c207 n90__i18__net4 vss 259.979e-18
c208 n85__i18__net4 vss 259.805e-18
c209 n82__i18__net4 vss 259.997e-18
c210 n75__i18__net4 vss 259.735e-18
c211 n70__i18__net4 vss 260.539e-18
c212 n65__i18__net4 vss 259.505e-18
c213 n61__i18__net4 vss 260.459e-18
c214 n55__i18__net4 vss 259.619e-18
c215 n50__i18__net4 vss 260.13e-18
c216 n47__i18__net4 vss 255.74e-18
c217 n42__i18__net4 vss 278.875e-18
c218 n39__i18__net4 vss 256.237e-18
c219 n36__i18__net4 vss 279.779e-18
c220 n33__i18__net4 vss 260.361e-18
c221 n30__i18__net4 vss 261.057e-18
c222 n27__i18__net4 vss 260.781e-18
c223 n24__i18__net4 vss 259.459e-18
c224 n21__i18__net4 vss 260.237e-18
c225 n18__i18__net4 vss 258.958e-18
c226 n15__i18__net4 vss 258.733e-18
c227 n12__i18__net4 vss 260.704e-18
c228 n9__i18__net4 vss 399.298e-18
c229 n6__i18__net4 vss 267.74e-18
c230 n3__i18__net4 vss 305.98e-18
c231 n472__i18__net5 vss 323.756e-18
c232 n465__i18__net5 vss 287.217e-18
c233 n460__i18__net5 vss 277.959e-18
c234 n455__i18__net5 vss 280.341e-18
c235 n452__i18__net5 vss 278.074e-18
c236 n445__i18__net5 vss 277.239e-18
c237 n442__i18__net5 vss 279.823e-18
c238 n437__i18__net5 vss 277.976e-18
c239 n430__i18__net5 vss 279.745e-18
c240 n425__i18__net5 vss 278.019e-18
c241 n421__i18__net5 vss 279.928e-18
c242 n415__i18__net5 vss 277.773e-18
c243 n410__i18__net5 vss 280.201e-18
c244 n407__i18__net5 vss 279.859e-18
c245 n400__i18__net5 vss 278.62e-18
c246 n397__i18__net5 vss 278.856e-18
c247 n392__i18__net5 vss 277.986e-18
c248 n387__i18__net5 vss 277.848e-18
c249 n380__i18__net5 vss 280.654e-18
c250 n377__i18__net5 vss 278.419e-18
c251 n370__i18__net5 vss 280.838e-18
c252 n367__i18__net5 vss 278.33e-18
c253 n362__i18__net5 vss 279.064e-18
c254 n357__i18__net5 vss 278.501e-18
c255 n350__i18__net5 vss 279.268e-18
c256 n347__i18__net5 vss 277.812e-18
c257 n340__i18__net5 vss 279.742e-18
c258 n337__i18__net5 vss 277.916e-18
c259 n330__i18__net5 vss 280.404e-18
c260 n327__i18__net5 vss 279.852e-18
c261 n322__i18__net5 vss 278.559e-18
c262 n315__i18__net5 vss 279.173e-18
c263 n312__i18__net5 vss 277.831e-18
c264 n305__i18__net5 vss 278.12e-18
c265 n300__i18__net5 vss 280.897e-18
c266 n295__i18__net5 vss 278.497e-18
c267 n290__i18__net5 vss 280.812e-18
c268 n285__i18__net5 vss 278.397e-18
c269 n280__i18__net5 vss 279.014e-18
c270 n277__i18__net5 vss 277.902e-18
c271 n270__i18__net5 vss 279.883e-18
c272 n267__i18__net5 vss 278.034e-18
c273 n260__i18__net5 vss 280.408e-18
c274 n255__i18__net5 vss 279.909e-18
c275 n252__i18__net5 vss 278.617e-18
c276 n247__i18__net5 vss 278.993e-18
c277 n242__i18__net5 vss 277.956e-18
c278 n237__i18__net5 vss 290.544e-18
c279 n230__i18__net5 vss 280.716e-18
c280 n225__i18__net5 vss 278.494e-18
c281 n220__i18__net5 vss 280.86e-18
c282 n216__i18__net5 vss 278.4e-18
c283 n210__i18__net5 vss 278.989e-18
c284 n205__i18__net5 vss 278.506e-18
c285 n201__i18__net5 vss 279.269e-18
c286 n195__i18__net5 vss 277.845e-18
c287 n190__i18__net5 vss 279.818e-18
c288 n187__i18__net5 vss 278.088e-18
c289 n181__i18__net5 vss 280.329e-18
c290 n175__i18__net5 vss 279.863e-18
c291 n172__i18__net5 vss 278.516e-18
c292 n166__i18__net5 vss 279.173e-18
c293 n162__i18__net5 vss 277.831e-18
c294 n155__i18__net5 vss 270.592e-18
c295 n150__i18__net5 vss 273.369e-18
c296 n145__i18__net5 vss 270.969e-18
c297 n140__i18__net5 vss 273.285e-18
c298 n137__i18__net5 vss 270.87e-18
c299 n131__i18__net5 vss 279.668e-18
c300 n125__i18__net5 vss 271.742e-18
c301 n122__i18__net5 vss 270.407e-18
c302 n117__i18__net5 vss 270.179e-18
c303 n112__i18__net5 vss 270.612e-18
c304 n105__i18__net5 vss 273.205e-18
c305 n102__i18__net5 vss 270.875e-18
c306 n97__i18__net5 vss 272.593e-18
c307 n92__i18__net5 vss 270.464e-18
c308 n87__i18__net5 vss 269.82e-18
c309 n80__i18__net5 vss 272.217e-18
c310 n75__i18__net5 vss 270.455e-18
c311 n70__i18__net5 vss 280.524e-18
c312 n65__i18__net5 vss 279.96e-18
c313 n62__i18__net5 vss 278.367e-18
c314 n55__i18__net5 vss 273.079e-18
c315 n52__i18__net5 vss 269.664e-18
c316 n45__i18__net5 vss 269.858e-18
c317 n42__i18__net5 vss 269.378e-18
c318 n39__i18__net5 vss 270.288e-18
c319 n36__i18__net5 vss 269.214e-18
c320 n33__i18__net5 vss 271.82e-18
c321 n30__i18__net5 vss 269.588e-18
c322 n27__i18__net5 vss 271.625e-18
c323 n24__i18__net5 vss 269.21e-18
c324 n21__i18__net5 vss 268.661e-18
c325 n18__i18__net5 vss 271.229e-18
c326 n15__i18__net5 vss 360.121e-18
c327 n12__i18__net5 vss 271.763e-18
c328 n9__i18__net5 vss 270.985e-18
c329 n6__i18__net5 vss 277.366e-18
c330 n3__i18__net5 vss 308.854e-18
c331 n6__net6 vss 21.7259e-18
c332 n8__net7 vss 15.6768e-18
c333 n7__net6 vss 14.7703e-18
c334 n8__net8 vss 14.7595e-18
c335 n10__net7 vss 20.4601e-18
c336 n9__net6 vss 18.5962e-18
c337 n10__net8 vss 18.6845e-18
c338 n10__r0 vss 29.7397e-18
c339 n8__r2 vss 26.3104e-18
c340 n13__serial_out vss 37.9869e-18
c341 n7__serial_out vss 24.0358e-18
c342 n11__net4 vss 26.3101e-18
c343 n6__net3 vss 26.3464e-18
c344 n4__i2__net77 vss 28.5156e-18
c345 n6__i1__net77 vss 30.3719e-18
c346 n4__i0__net77 vss 31.65e-18
c347 n5__i1__net76 vss 22.5995e-18
c348 n7__i2__net76 vss 23.587e-18
c349 n6__i1__net76 vss 26.3822e-18
c350 n7__i0__net76 vss 26.0801e-18
c351 n15__reset_b vss 17.5032e-18
c352 n17__reset_b vss 16.821e-18
c353 n19__reset_b vss 16.6115e-18
c354 n3__i2__net77 vss 31.3451e-18
c355 n2__i1__net77 vss 30.8354e-18
c356 n3__i0__net77 vss 30.4388e-18
c357 n8__i13__net7 vss 25.7384e-18
c358 n9__i13__net18 vss 19.8659e-18
c359 n26__ck_b vss 16.6379e-18
c360 n28__ck_b vss 17.9829e-18
c361 n30__ck_b vss 17.8988e-18
c362 n8__i13__net18 vss 22.74e-18
c363 n5__i1__net74 vss 26.8843e-18
c364 n7__i2__net74 vss 23.4481e-18
c365 n6__i1__net74 vss 26.2686e-18
c366 n7__i0__net74 vss 26.1803e-18
c367 n4__i13__i20__net1 vss 27.6354e-18
c368 n4__i13__net18 vss 44.5605e-18
c369 n4__i13__net7 vss 33.9724e-18
c370 n3__i2__net75 vss 30.6867e-18
c371 n2__i1__net75 vss 32.9971e-18
c372 n3__i0__net75 vss 31.2141e-18
c373 n17__ck_buff vss 19.3261e-18
c374 n19__ck_buff vss 17.747e-18
c375 n21__ck_buff vss 17.7148e-18
c376 n8__i13__net11 vss 23.4951e-18
c377 n5__i13__net12 vss 21.4128e-18
c378 n9__i13__net1 vss 19.7631e-18
c379 n9__i13__net2 vss 19.5709e-18
c380 n4__i1__net1 vss 30.8249e-18
c381 n8__i13__net1 vss 22.4259e-18
c382 n5__i13__net2 vss 22.4976e-18
c383 n4__i13__i19__net1 vss 26.4835e-18
c384 n20__shift vss 30.685e-18
c385 n22__shift vss 29.003e-18
c386 n24__shift vss 28.2864e-18
c387 n4__i13__net1 vss 44.0725e-18
c388 n4__i13__net11 vss 34.3888e-18
c389 n8__shift vss 31.4212e-18
c390 n9__shift vss 30.9343e-18
c391 n10__ck4 vss 22.1756e-18
c392 n15__ck4 vss 30.6848e-18
c393 n8__i13__a3 vss 23.2643e-18
c394 n5__i13__a1 vss 23.1745e-18
c395 n3__net14 vss 26.8425e-18
c396 n6__i9__net1 vss 16.034e-18
c397 n13__i13__a2 vss 19.7442e-18
c398 n13__i13__a0 vss 19.712e-18
c399 n5__net14 vss 17.144e-18
c400 n7__net14 vss 22.9061e-18
c401 n8__i13__a2 vss 22.9718e-18
c402 n5__i13__a0 vss 23.0273e-18
c403 n3__net13 vss 23.785e-18
c404 n5__net13 vss 16.439e-18
c405 n58__reset vss 24.9569e-18
c406 n4__i9__i4__net4 vss 32.2454e-18
c407 n7__net13 vss 26.902e-18
c408 n4__i13__i17__net1 vss 27.467e-18
c409 n4__i13__a2 vss 44.6173e-18
c410 n53__reset vss 26.7449e-18
c411 n29__ck vss 24.0293e-18
c412 n7__i9__i4__net5 vss 28.116e-18
c413 n4__i13__a3 vss 33.6165e-18
c414 n6__net10 vss 20.6705e-18
c415 n8__net10 vss 16.1015e-18
c416 n5__net10 vss 19.7542e-18
c417 n3__i9__i4__net4 vss 31.201e-18
c418 n4__y_out_3 vss 24.315e-18
c419 n5__net12 vss 22.7834e-18
c420 n4__ck_b vss 16.9192e-18
c421 n7__net12 vss 17.3076e-18
c422 n10__x_out_3 vss 19.6299e-18
c423 n10__x_out_1 vss 19.6677e-18
c424 n9__net12 vss 25.8056e-18
c425 n24__ck vss 28.1938e-18
c426 n7__i9__i4__net1 vss 25.6822e-18
c427 n9__x_out_3 vss 20.2628e-18
c428 n6__x_out_1 vss 20.1672e-18
c429 n6__net9 vss 20.1934e-18
c430 n8__net9 vss 14.4101e-18
c431 n5__net9 vss 18.5501e-18
c432 n4__y_out_2 vss 22.2699e-18
c433 n6__x_out_0 vss 21.6727e-18
c434 n3__i9__i4__net2 vss 31.9983e-18
c435 n10__x_out_2 vss 19.4809e-18
c436 n5__y_out_0 vss 19.5406e-18
c437 n5__net11 vss 23.4488e-18
c438 n2__ck_buff vss 20.4432e-18
c439 n7__net11 vss 19.6282e-18
c440 n9__net11 vss 23.4803e-18
c441 n9__x_out_2 vss 20.4211e-18
c442 n15__i14__net7 vss 22.1272e-18
c443 n5__i14__net11 vss 27.2098e-18
c444 n4__i14__x_out_b_1 vss 27.7594e-18
c445 n4__i14__y_out_b_1 vss 28.6974e-18
c446 n16__i14__net7 vss 17.7146e-18
c447 n17__i14__net11 vss 18.9796e-18
c448 n18__i14__net7 vss 18.6289e-18
c449 n19__i14__net11 vss 18.8816e-18
c450 n6__i14__i11__net4 vss 30.0395e-18
c451 n4__i14__i14__net4 vss 31.4048e-18
c452 n6__i14__i15__net4 vss 30.0628e-18
c453 n4__i14__i12__net4 vss 31.4291e-18
c454 n20__i14__net7 vss 18.9168e-18
c455 n21__i14__net11 vss 19.3893e-18
c456 n22__i14__net7 vss 18.5382e-18
c457 n23__i14__net11 vss 18.722e-18
c458 n5__i14__i11__net5 vss 23.0224e-18
c459 n5__i14__i15__net5 vss 23.0773e-18
c460 n14__i14__net7 vss 24.5584e-18
c461 n24__i14__net11 vss 24.3573e-18
c462 n6__i14__i11__net5 vss 26.3916e-18
c463 n7__i14__i14__net5 vss 26.3689e-18
c464 n6__i14__i15__net5 vss 26.3916e-18
c465 n7__i14__i12__net5 vss 26.3689e-18
c466 n29__i14__net4 vss 25.6151e-18
c467 n4__i14__net11 vss 30.4256e-18
c468 n21__i14__net4 vss 16.1491e-18
c469 n23__i14__net4 vss 16.1491e-18
c470 n25__i14__net4 vss 16.1491e-18
c471 n27__i14__net4 vss 16.1491e-18
c472 n41__i14__net4 vss 17.8866e-18
c473 n43__i14__net4 vss 14.9656e-18
c474 n4__i14__net7 vss 29.1935e-18
c475 n2__i14__i11__net4 vss 30.2474e-18
c476 n3__i14__i14__net4 vss 29.744e-18
c477 n2__i14__i15__net4 vss 30.2523e-18
c478 n3__i14__i12__net4 vss 29.744e-18
c479 n45__i14__net4 vss 20.5345e-18
c480 n47__i14__net4 vss 15.0491e-18
c481 n48__i14__net4 vss 25.4854e-18
c482 n50__i14__net9 vss 16.6823e-18
c483 n52__i14__net9 vss 16.6235e-18
c484 n54__i14__net9 vss 16.6823e-18
c485 n56__i14__net9 vss 16.6235e-18
c486 n36__reset vss 20.9185e-18
c487 n6__i14__i17__net11 vss 37.6501e-18
c488 n37__reset vss 19.2009e-18
c489 n5__i14__i11__net1 vss 26.819e-18
c490 n5__i14__i15__net1 vss 26.819e-18
c491 n15__i14__i17__net8 vss 40.9128e-18
c492 n39__reset vss 18.8696e-18
c493 n6__i14__i11__net1 vss 24.7933e-18
c494 n7__i14__i14__net1 vss 24.7688e-18
c495 n6__i14__i15__net1 vss 24.7933e-18
c496 n7__i14__i12__net1 vss 24.7677e-18
c497 n41__reset vss 15.8447e-18
c498 n43__reset vss 17.3733e-18
c499 n5__i14__i17__net10 vss 28.0174e-18
c500 n35__reset vss 21.7972e-18
c501 n5__i14__i17__net9 vss 29.0962e-18
c502 n4__i14__i17__net9 vss 27.8945e-18
c503 n2__i14__i17__net11 vss 50.4804e-18
c504 n2__i14__i11__net2 vss 28.9261e-18
c505 n3__i14__i14__net2 vss 28.2135e-18
c506 n2__i14__i15__net2 vss 28.9261e-18
c507 n3__i14__i12__net2 vss 28.2135e-18
c508 n4__i14__i17__net10 vss 30.6943e-18
c509 n10__i14__i17__net8 vss 28.7659e-18
c510 n30__i14__net10 vss 17.3312e-18
c511 n32__i14__net10 vss 17.3312e-18
c512 n34__i14__net10 vss 17.3312e-18
c513 n36__i14__net10 vss 17.3312e-18
c514 n17__i14__i17__net1 vss 26.8105e-18
c515 n6__i14__i17__net8 vss 25.5687e-18
c516 n6__i14__i17__i2__net4 vss 29.446e-18
c517 n4__i14__i17__i3__net4 vss 32.321e-18
c518 n4__i14__y_out_b_3 vss 30.4966e-18
c519 n4__i14__x_out_b_2 vss 30.4966e-18
c520 n5__i14__i17__i2__net5 vss 22.0518e-18
c521 n6__i14__i13__net4 vss 29.531e-18
c522 n4__i14__i16__net4 vss 30.9417e-18
c523 n6__i14__i10__net4 vss 29.5733e-18
c524 n4__i14__i9__net4 vss 30.9417e-18
c525 n6__i14__i17__i2__net5 vss 26.929e-18
c526 n7__i14__i17__i3__net5 vss 25.5608e-18
c527 n5__i14__i13__net5 vss 22.6899e-18
c528 n5__i14__i10__net5 vss 22.6899e-18
c529 n3__i14__i17__net6 vss 18.0505e-18
c530 n6__i14__i13__net5 vss 26.4304e-18
c531 n7__i14__i16__net5 vss 26.4079e-18
c532 n6__i14__i10__net5 vss 26.4304e-18
c533 n7__i14__i9__net5 vss 26.4079e-18
c534 n2__i14__i17__i2__net4 vss 30.5959e-18
c535 n3__i14__i17__i3__net4 vss 30.862e-18
c536 n3__i14__net4 vss 16.5107e-18
c537 n5__i14__net4 vss 16.5107e-18
c538 n7__i14__net4 vss 16.5107e-18
c539 n2__i14__i13__net4 vss 31.2785e-18
c540 n3__i14__i16__net4 vss 32.2898e-18
c541 n2__i14__i10__net4 vss 32.329e-18
c542 n3__i14__i9__net4 vss 32.2929e-18
c543 n4__i14__i17__net3 vss 19.1434e-18
c544 n4__i14__i17__net1 vss 19.0215e-18
c545 n5__i14__i17__i2__net1 vss 26.3223e-18
c546 n10__i14__net9 vss 16.9789e-18
c547 n12__i14__net9 vss 16.92e-18
c548 n14__i14__net9 vss 16.953e-18
c549 n16__i14__net9 vss 16.8941e-18
c550 n6__i14__i17__i2__net1 vss 24.8206e-18
c551 n7__i14__i17__i3__net1 vss 25.019e-18
c552 n5__i14__i13__net1 vss 26.2939e-18
c553 n5__i14__i10__net1 vss 26.2939e-18
c554 n6__i14__i13__net1 vss 25.5452e-18
c555 n7__i14__i16__net1 vss 25.5479e-18
c556 n6__i14__i10__net1 vss 25.5725e-18
c557 n7__i14__i9__net1 vss 25.5479e-18
c558 n2__i14__i17__i2__net2 vss 28.8734e-18
c559 n3__i14__i17__i3__net2 vss 28.3945e-18
c560 n2__i14__i13__net2 vss 31.2049e-18
c561 n3__i14__i16__net2 vss 30.5513e-18
c562 n2__i14__i10__net2 vss 31.2468e-18
c563 n3__i14__i9__net2 vss 30.4935e-18
c564 n5__ck vss 16.9411e-18
c565 n2__i14__i17__net7 vss 19.2894e-18
c566 n3__ck vss 20.0886e-18
c567 n1__reset vss 39.0429e-18
c568 n2__i14__net10 vss 17.4906e-18
c569 n4__i14__net10 vss 17.3679e-18
c570 n6__i14__net10 vss 17.4906e-18
c571 n8__i14__net10 vss 17.3679e-18
c572 n4__serial_out_b_high vss 34.9644e-18
c573 n6__i18__net1 vss 94.5229e-18
c574 n6__i12__bcore_bar vss 24.9238e-18
c575 n4__i12__bcore_bar vss 19.796e-18
c576 n9__i18__net2 vss 120.575e-18
c577 n2__i12__bcore_bar vss 24.7604e-18
c578 n11__i18__net2 vss 120.412e-18
c579 n12__i18__net2 vss 151.333e-18
c580 n6__serial_out vss 25.5124e-18
c581 n4__serial_out vss 19.9498e-18
c582 n2__serial_out vss 25.7759e-18
c583 n28__i18__net3 vss 201.604e-18
c584 n25__i18__net3 vss 163.292e-18
c585 n22__i18__net3 vss 163.861e-18
c586 n19__i18__net3 vss 164.265e-18
c587 n16__i18__net3 vss 164.324e-18
c588 n13__i18__net3 vss 164.224e-18
c589 n10__i18__net3 vss 163.526e-18
c590 n7__i18__net3 vss 164.124e-18
c591 n4__i18__net3 vss 168.529e-18
c592 n120__i18__net4 vss 246.967e-18
c593 n113__i18__net4 vss 199.451e-18
c594 n110__i18__net4 vss 195.584e-18
c595 n103__i18__net4 vss 194.808e-18
c596 n100__i18__net4 vss 190.226e-18
c597 n95__i18__net4 vss 195.806e-18
c598 n88__i18__net4 vss 190.344e-18
c599 n83__i18__net4 vss 196.313e-18
c600 n80__i18__net4 vss 196.137e-18
c601 n73__i18__net4 vss 203.622e-18
c602 n68__i18__net4 vss 191.099e-18
c603 n63__i18__net4 vss 195.982e-18
c604 n59__i18__net4 vss 196.177e-18
c605 n53__i18__net4 vss 195.706e-18
c606 n48__i18__net4 vss 193.047e-18
c607 n45__i18__net4 vss 190.777e-18
c608 n40__i18__net4 vss 204.367e-18
c609 n37__i18__net4 vss 192.339e-18
c610 n34__i18__net4 vss 205.562e-18
c611 n31__i18__net4 vss 196.401e-18
c612 n28__i18__net4 vss 190.565e-18
c613 n25__i18__net4 vss 196.829e-18
c614 n22__i18__net4 vss 195.193e-18
c615 n19__i18__net4 vss 196.706e-18
c616 n16__i18__net4 vss 195.451e-18
c617 n13__i18__net4 vss 194.07e-18
c618 n10__i18__net4 vss 196.725e-18
c619 n7__i18__net4 vss 213.263e-18
c620 n4__i18__net4 vss 200.378e-18
c621 n470__i18__net5 vss 246.4e-18
c622 n463__i18__net5 vss 218.318e-18
c623 n458__i18__net5 vss 200.679e-18
c624 n453__i18__net5 vss 209.875e-18
c625 n450__i18__net5 vss 212.044e-18
c626 n443__i18__net5 vss 207.86e-18
c627 n440__i18__net5 vss 212.07e-18
c628 n435__i18__net5 vss 259.097e-18
c629 n428__i18__net5 vss 213.494e-18
c630 n423__i18__net5 vss 206.842e-18
c631 n419__i18__net5 vss 211.834e-18
c632 n413__i18__net5 vss 211.585e-18
c633 n408__i18__net5 vss 208.696e-18
c634 n405__i18__net5 vss 211.678e-18
c635 n398__i18__net5 vss 207.158e-18
c636 n395__i18__net5 vss 209.718e-18
c637 n390__i18__net5 vss 209.948e-18
c638 n385__i18__net5 vss 211.616e-18
c639 n378__i18__net5 vss 209.399e-18
c640 n375__i18__net5 vss 212.334e-18
c641 n368__i18__net5 vss 215.142e-18
c642 n365__i18__net5 vss 209.133e-18
c643 n360__i18__net5 vss 207.992e-18
c644 n355__i18__net5 vss 213.419e-18
c645 n348__i18__net5 vss 213.233e-18
c646 n345__i18__net5 vss 211.359e-18
c647 n338__i18__net5 vss 213.387e-18
c648 n335__i18__net5 vss 211.603e-18
c649 n328__i18__net5 vss 213.88e-18
c650 n325__i18__net5 vss 213.339e-18
c651 n320__i18__net5 vss 212.118e-18
c652 n313__i18__net5 vss 212.654e-18
c653 n310__i18__net5 vss 211.369e-18
c654 n303__i18__net5 vss 211.617e-18
c655 n298__i18__net5 vss 214.309e-18
c656 n293__i18__net5 vss 212.053e-18
c657 n288__i18__net5 vss 214.269e-18
c658 n283__i18__net5 vss 211.851e-18
c659 n278__i18__net5 vss 212.468e-18
c660 n275__i18__net5 vss 211.427e-18
c661 n268__i18__net5 vss 213.373e-18
c662 n265__i18__net5 vss 211.577e-18
c663 n258__i18__net5 vss 213.896e-18
c664 n253__i18__net5 vss 213.416e-18
c665 n250__i18__net5 vss 212.142e-18
c666 n245__i18__net5 vss 212.514e-18
c667 n240__i18__net5 vss 211.596e-18
c668 n235__i18__net5 vss 211.618e-18
c669 n228__i18__net5 vss 214.171e-18
c670 n223__i18__net5 vss 212.018e-18
c671 n218__i18__net5 vss 214.327e-18
c672 n214__i18__net5 vss 211.866e-18
c673 n208__i18__net5 vss 212.443e-18
c674 n203__i18__net5 vss 212.038e-18
c675 n199__i18__net5 vss 212.683e-18
c676 n193__i18__net5 vss 211.443e-18
c677 n188__i18__net5 vss 213.326e-18
c678 n185__i18__net5 vss 211.631e-18
c679 n179__i18__net5 vss 213.817e-18
c680 n173__i18__net5 vss 213.361e-18
c681 n170__i18__net5 vss 212.116e-18
c682 n164__i18__net5 vss 212.654e-18
c683 n160__i18__net5 vss 211.333e-18
c684 n153__i18__net5 vss 211.617e-18
c685 n148__i18__net5 vss 214.309e-18
c686 n143__i18__net5 vss 212.013e-18
c687 n138__i18__net5 vss 214.354e-18
c688 n135__i18__net5 vss 211.942e-18
c689 n129__i18__net5 vss 226.891e-18
c690 n123__i18__net5 vss 212.784e-18
c691 n120__i18__net5 vss 211.535e-18
c692 n115__i18__net5 vss 211.539e-18
c693 n110__i18__net5 vss 210.537e-18
c694 n103__i18__net5 vss 214.21e-18
c695 n100__i18__net5 vss 211.86e-18
c696 n95__i18__net5 vss 213.741e-18
c697 n90__i18__net5 vss 211.605e-18
c698 n85__i18__net5 vss 210.871e-18
c699 n78__i18__net5 vss 213.2e-18
c700 n73__i18__net5 vss 211.507e-18
c701 n68__i18__net5 vss 214.027e-18
c702 n63__i18__net5 vss 213.474e-18
c703 n60__i18__net5 vss 211.903e-18
c704 n53__i18__net5 vss 212.28e-18
c705 n50__i18__net5 vss 207.468e-18
c706 n43__i18__net5 vss 207.593e-18
c707 n40__i18__net5 vss 207.296e-18
c708 n37__i18__net5 vss 208.134e-18
c709 n34__i18__net5 vss 207.043e-18
c710 n31__i18__net5 vss 209.874e-18
c711 n28__i18__net5 vss 207.552e-18
c712 n25__i18__net5 vss 209.512e-18
c713 n22__i18__net5 vss 207.103e-18
c714 n19__i18__net5 vss 206.551e-18
c715 n16__i18__net5 vss 209.051e-18
c716 n13__i18__net5 vss 207.159e-18
c717 n10__i18__net5 vss 209.757e-18
c718 n7__i18__net5 vss 208.901e-18
c719 n4__i18__net5 vss 213.233e-18
c720 n6__net7 vss 18.9555e-18
c721 n6__net8 vss 18.835e-18
c722 n7__net7 vss 12.7425e-18
c723 n8__net6 vss 13.0373e-18
c724 n7__net8 vss 12.8926e-18
c725 n9__net7 vss 16.5958e-18
c726 n10__net6 vss 16.8433e-18
c727 n9__net8 vss 18.0045e-18
c728 n13__r0 vss 23.8431e-18
c729 n5__r2 vss 23.8119e-18
c730 n4__r1 vss 25.0112e-18
c731 n11__serial_out vss 23.5754e-18
c732 n10__serial_out vss 20.8736e-18
c733 n8__net4 vss 20.5368e-18
c734 n9__net3 vss 19.4485e-18
c735 n6__i2__net77 vss 23.9163e-18
c736 n4__i1__net77 vss 24.2223e-18
c737 n6__i0__net77 vss 21.9733e-18
c738 n5__i2__net76 vss 17.6939e-18
c739 n5__i0__net76 vss 16.5918e-18
c740 n6__i2__net76 vss 22.2699e-18
c741 n7__i1__net76 vss 20.6176e-18
c742 n6__i0__net76 vss 20.3798e-18
c743 n2__i2__net77 vss 77.2528e-18
c744 n3__i1__net77 vss 72.4297e-18
c745 n2__i0__net77 vss 74.5151e-18
c746 n5__i13__net7 vss 19.8472e-18
c747 n29__ck_buff vss 23.4441e-18
c748 n31__ck_buff vss 22.9522e-18
c749 n33__ck_buff vss 22.9114e-18
c750 n5__i13__net18 vss 22.6068e-18
c751 n5__i2__net74 vss 19.7306e-18
c752 n5__i0__net74 vss 19.6883e-18
c753 n6__i2__net74 vss 21.2597e-18
c754 n7__i1__net74 vss 21.041e-18
c755 n6__i0__net74 vss 20.2427e-18
c756 n3__i13__net3 vss 26.8486e-18
c757 n21__reset_buff vss 23.0607e-18
c758 n23__reset_buff vss 22.6016e-18
c759 n25__reset_buff vss 25.8464e-18
c760 n4__i13__net23 vss 25.2829e-18
c761 n2__i2__net75 vss 76.7775e-18
c762 n3__i1__net75 vss 72.6882e-18
c763 n2__i0__net75 vss 79.3923e-18
c764 n4__i13__net17 vss 37.5384e-18
c765 n20__ck_b vss 20.5971e-18
c766 n22__ck_b vss 20.6807e-18
c767 n24__ck_b vss 24.0067e-18
c768 n5__i13__net11 vss 22.0186e-18
c769 n8__i13__net12 vss 20.404e-18
c770 n4__i2__net1 vss 23.8054e-18
c771 n4__i0__net1 vss 25.6771e-18
c772 n5__i13__net1 vss 23.4544e-18
c773 n8__i13__net2 vss 25.1079e-18
c774 n4__i13__i18__net1 vss 22.3134e-18
c775 n3__i2__net79 vss 24.7988e-18
c776 n3__i1__net79 vss 26.487e-18
c777 n3__i0__net79 vss 24.9697e-18
c778 n4__i13__net2 vss 30.9471e-18
c779 n13__shift vss 28.6265e-18
c780 n15__shift vss 28.6378e-18
c781 n17__shift vss 29.9074e-18
c782 n4__i13__net12 vss 44.6243e-18
c783 n4__shift vss 16.3964e-18
c784 n5__shift vss 16.6952e-18
c785 n12__shift vss 20.8009e-18
c786 n13__ck4 vss 25.6773e-18
c787 n14__ck4 vss 31.6317e-18
c788 n5__i13__a3 vss 21.5104e-18
c789 n8__i13__a1 vss 19.681e-18
c790 n4__i9__net1 vss 29.5295e-18
c791 n5__i9__net1 vss 22.8796e-18
c792 n8__net14 vss 12.338e-18
c793 n10__net14 vss 18.1111e-18
c794 n5__i13__a2 vss 24.9754e-18
c795 n8__i13__a0 vss 23.1981e-18
c796 n4__i9__net2 vss 22.6048e-18
c797 n8__net13 vss 11.1894e-18
c798 n55__reset vss 20.5564e-18
c799 n6__i9__i4__net4 vss 20.3419e-18
c800 n10__net13 vss 17.5575e-18
c801 n4__i13__i16__net1 vss 24.6348e-18
c802 n5__i9__i4__net5 vss 16.8267e-18
c803 n4__i13__a0 vss 34.3965e-18
c804 n54__reset vss 22.5257e-18
c805 n26__ck vss 23.836e-18
c806 n6__i9__i4__net5 vss 19.2595e-18
c807 n4__i13__a1 vss 40.9855e-18
c808 n7__net10 vss 17.3838e-18
c809 n2__i9__i4__net4 vss 75.2536e-18
c810 n9__net10 vss 13.5706e-18
c811 n10__net10 vss 16.3741e-18
c812 n4__y_out_1 vss 18.3043e-18
c813 n6__net12 vss 19.9996e-18
c814 n4__ck_buff vss 24.4505e-18
c815 n8__net12 vss 11.5919e-18
c816 n10__net12 vss 16.733e-18
c817 n5__i9__i4__net1 vss 19.4973e-18
c818 n25__ck vss 27.0715e-18
c819 n6__i9__i4__net1 vss 22.0225e-18
c820 n6__x_out_3 vss 20.7348e-18
c821 n9__x_out_1 vss 22.5276e-18
c822 n2__reset_buff vss 24.8792e-18
c823 n7__net9 vss 18.8002e-18
c824 n2__i9__i4__net2 vss 76.1202e-18
c825 n9__net9 vss 14.2491e-18
c826 n10__net9 vss 17.3294e-18
c827 n9__x_out_0 vss 17.9591e-18
c828 n6__net11 vss 17.2814e-18
c829 n2__ck_b vss 24.4814e-18
c830 n8__net11 vss 12.2146e-18
c831 n10__net11 vss 17.9378e-18
c832 n6__x_out_2 vss 22.2666e-18
c833 n4__y_out_0 vss 20.0412e-18
c834 n5__i14__net7 vss 16.6515e-18
c835 n15__i14__net11 vss 17.7757e-18
c836 n4__i14__y_out_b_2 vss 21.9734e-18
c837 n4__i14__x_out_b_0 vss 21.1594e-18
c838 n17__i14__net7 vss 12.0737e-18
c839 n16__i14__net11 vss 13.6268e-18
c840 n19__i14__net7 vss 11.8838e-18
c841 n18__i14__net11 vss 12.7931e-18
c842 n4__i14__i11__net4 vss 27.0659e-18
c843 n6__i14__i14__net4 vss 23.4914e-18
c844 n4__i14__i15__net4 vss 25.0942e-18
c845 n6__i14__i12__net4 vss 24.6787e-18
c846 n21__i14__net7 vss 11.8759e-18
c847 n20__i14__net11 vss 12.6114e-18
c848 n23__i14__net7 vss 11.8694e-18
c849 n22__i14__net11 vss 11.9394e-18
c850 n5__i14__i14__net5 vss 17.1594e-18
c851 n5__i14__i12__net5 vss 15.6966e-18
c852 n24__i14__net7 vss 17.3013e-18
c853 n14__i14__net11 vss 19.334e-18
c854 n7__i14__i11__net5 vss 21.708e-18
c855 n6__i14__i14__net5 vss 22.5411e-18
c856 n7__i14__i15__net5 vss 22.515e-18
c857 n6__i14__i12__net5 vss 19.3042e-18
c858 n39__i14__net4 vss 15.914e-18
c859 n40__i14__net4 vss 14.7545e-18
c860 n3__i14__i11__net4 vss 71.482e-18
c861 n2__i14__i14__net4 vss 71.8362e-18
c862 n3__i14__i15__net4 vss 71.2793e-18
c863 n2__i14__i12__net4 vss 71.1217e-18
c864 n42__i14__net4 vss 15.5034e-18
c865 n44__i14__net4 vss 16.4291e-18
c866 n46__i14__net4 vss 12.0074e-18
c867 n38__i14__net4 vss 18.1755e-18
c868 n58__i14__net10 vss 25.6223e-18
c869 n60__i14__net10 vss 22.6563e-18
c870 n62__i14__net10 vss 22.5171e-18
c871 n64__i14__net10 vss 24.4074e-18
c872 n26__reset vss 15.9275e-18
c873 n14__i14__i17__net8 vss 52.1514e-18
c874 n38__reset vss 11.9507e-18
c875 n5__i14__i14__net1 vss 19.0524e-18
c876 n5__i14__i12__net1 vss 19.8459e-18
c877 n4__i14__i17__net11 vss 26.4631e-18
c878 n40__reset vss 11.7395e-18
c879 n7__i14__i11__net1 vss 19.6348e-18
c880 n6__i14__i14__net1 vss 20.6473e-18
c881 n7__i14__i15__net1 vss 20.654e-18
c882 n6__i14__i12__net1 vss 21.2323e-18
c883 n42__reset vss 11.4907e-18
c884 n44__reset vss 11.7229e-18
c885 n7__i14__i17__net10 vss 25.3019e-18
c886 n30__i14__net3 vss 23.7642e-18
c887 n32__i14__net3 vss 22.1025e-18
c888 n34__i14__net3 vss 21.9763e-18
c889 n36__i14__net3 vss 23.8439e-18
c890 n45__reset vss 16.7636e-18
c891 n7__i14__i17__net9 vss 22.004e-18
c892 n3__i14__i11__net2 vss 71.8751e-18
c893 n2__i14__i14__net2 vss 72.8249e-18
c894 n3__i14__i15__net2 vss 72.6954e-18
c895 n2__i14__i12__net2 vss 73.2492e-18
c896 n13__i14__i17__net8 vss 26.3888e-18
c897 n3__i14__i17__net11 vss 47.3384e-18
c898 n34__i14__net9 vss 25.1404e-18
c899 n36__i14__net9 vss 21.7273e-18
c900 n38__i14__net9 vss 21.5649e-18
c901 n40__i14__net9 vss 24.4437e-18
c902 n14__i14__i17__net1 vss 20.0186e-18
c903 n9__i14__i17__net8 vss 23.2939e-18
c904 n4__i14__i17__i2__net4 vss 22.3441e-18
c905 n6__i14__i17__i3__net4 vss 24.9339e-18
c906 n4__i14__y_out_b_0 vss 21.8776e-18
c907 n4__i14__x_out_b_3 vss 20.2803e-18
c908 n5__i14__i17__i3__net5 vss 19.2255e-18
c909 n4__i14__i13__net4 vss 26.5892e-18
c910 n6__i14__i16__net4 vss 23.4371e-18
c911 n4__i14__i10__net4 vss 24.9679e-18
c912 n6__i14__i9__net4 vss 26.0372e-18
c913 n7__i14__i17__i2__net5 vss 20.5096e-18
c914 n6__i14__i17__i3__net5 vss 21.7577e-18
c915 n5__i14__i16__net5 vss 17.3213e-18
c916 n5__i14__i9__net5 vss 15.8188e-18
c917 n7__i14__i13__net5 vss 22.6196e-18
c918 n6__i14__i16__net5 vss 21.6953e-18
c919 n7__i14__i10__net5 vss 21.6691e-18
c920 n6__i14__i9__net5 vss 24.2706e-18
c921 n3__i14__i17__i2__net4 vss 69.7817e-18
c922 n2__i14__i17__i3__net4 vss 75.1516e-18
c923 n3__i14__i13__net4 vss 72.9357e-18
c924 n2__i14__i16__net4 vss 75.0074e-18
c925 n3__i14__i10__net4 vss 74.9152e-18
c926 n2__i14__i9__net4 vss 77.517e-18
c927 n7__ck vss 24.6101e-18
c928 n4__i14__i17__net7 vss 24.4821e-18
c929 n5__i14__i17__i3__net1 vss 20.4802e-18
c930 n10__i14__net10 vss 23.8708e-18
c931 n12__i14__net10 vss 23.3407e-18
c932 n14__i14__net10 vss 23.2074e-18
c933 n16__i14__net10 vss 25.7291e-18
c934 n7__i14__i17__i2__net1 vss 18.7469e-18
c935 n6__i14__i17__i3__net1 vss 19.3631e-18
c936 n5__i14__i16__net1 vss 19.6178e-18
c937 n5__i14__i9__net1 vss 18.1578e-18
c938 n5__reset vss 23.5444e-18
c939 n7__reset vss 23.0364e-18
c940 n7__i14__i13__net1 vss 23.4342e-18
c941 n6__i14__i16__net1 vss 20.7895e-18
c942 n7__i14__i10__net1 vss 20.7939e-18
c943 n6__i14__i9__net1 vss 21.4515e-18
c944 n3__i14__i17__i2__net2 vss 67.627e-18
c945 n2__i14__i17__i3__net2 vss 77.1314e-18
c946 n2__i14__net3 vss 23.7786e-18
c947 n4__i14__net3 vss 22.1992e-18
c948 n6__i14__net3 vss 22.073e-18
c949 n8__i14__net3 vss 24.2272e-18
c950 n3__i14__i13__net2 vss 76.7808e-18
c951 n2__i14__i16__net2 vss 80.5357e-18
c952 n3__i14__i10__net2 vss 80.4061e-18
c953 n2__i14__i9__net2 vss 87.4024e-18
c954 n2__i14__i17__net3 vss 24.9157e-18
c955 n2__i14__i17__net1 vss 25.8537e-18
c956 n1__ck vss 36.0982e-18
c957 n3__reset vss 26.3544e-18
c958 n2__i14__net9 vss 24.7338e-18
c959 n4__i14__net9 vss 25.2594e-18
c960 n6__i14__net9 vss 25.2594e-18
c961 n8__i14__net9 vss 28.0833e-18
c962 n2__serial_out_b_high_buff vss 68.3174e-18
c963 n3__serial_out_b_high vss 113.2e-18
c964 n5__net7 vss 69.4047e-18
c965 n5__net6 vss 70.847e-18
c966 n5__net8 vss 68.3271e-18
c967 n12__serial_out vss 41.646e-18
c968 n2__i18__net1 vss 92.6639e-18
c969 n12__r0 vss 49.138e-18
c970 n7__r2 vss 47.0008e-18
c971 n3__r1 vss 57.2407e-18
c972 n5__i12__bcore_bar vss 194.939e-18
c973 n2__i18__net2 vss 95.7141e-18
c974 n3__i12__bcore_bar vss 155.966e-18
c975 n9__serial_out vss 60.0703e-18
c976 n10__net4 vss 59.7531e-18
c977 n8__net3 vss 58.7364e-18
c978 n5__i2__net77 vss 20.8696e-18
c979 n5__i1__net77 vss 20.821e-18
c980 n5__i0__net77 vss 20.5869e-18
c981 n5__serial_out vss 262.46e-18
c982 n4__i2__net76 vss 83.7286e-18
c983 n4__i1__net76 vss 83.9569e-18
c984 n4__i0__net76 vss 81.3313e-18
c985 n3__serial_out vss 97.2428e-18
c986 n16__reset_b vss 46.3282e-18
c987 n18__reset_b vss 45.4204e-18
c988 n20__reset_b vss 44.945e-18
c989 n1__serial_out vss 105.241e-18
c990 n29__i18__net3 vss 18.394e-18
c991 n7__i13__net7 vss 99.2826e-18
c992 n26__i18__net3 vss 10.3882e-18
c993 n2__i13__i20__i4__net2 vss 22.4942e-18
c994 n25__ck_b vss 25.8437e-18
c995 n28__ck_buff vss 30.9087e-18
c996 n30__ck_buff vss 30.8359e-18
c997 n27__ck_b vss 26.3386e-18
c998 n29__ck_b vss 26.1879e-18
c999 n32__ck_buff vss 31.0735e-18
c1000 n10__i13__net18 vss 41.0703e-18
c1001 n23__i18__net3 vss 15.2412e-18
c1002 n20__i18__net3 vss 15.1974e-18
c1003 n7__i13__net18 vss 10.7429e-18
c1004 n4__i2__net74 vss 86.8615e-18
c1005 n4__i1__net74 vss 87.8089e-18
c1006 n4__i0__net74 vss 91.2651e-18
c1007 n17__i18__net3 vss 15.1974e-18
c1008 n2__i13__net3 vss 72.9027e-18
c1009 n3__i13__i20__net1 vss 53.2916e-18
c1010 n20__reset_buff vss 23.2865e-18
c1011 n22__reset_buff vss 23.2701e-18
c1012 n24__reset_buff vss 23.9757e-18
c1013 n14__i18__net3 vss 15.2169e-18
c1014 n3__i13__net23 vss 21.1504e-18
c1015 n3__i13__net18 vss 24.2767e-18
c1016 n11__i18__net3 vss 15.2169e-18
c1017 n3__i13__net17 vss 12.7457e-18
c1018 n3__i13__net7 vss 13.9608e-18
c1019 n8__i18__net3 vss 15.2169e-18
c1020 n5__i18__net3 vss 14.983e-18
c1021 n16__ck_buff vss 27.5069e-18
c1022 n19__ck_b vss 29.4679e-18
c1023 n21__ck_b vss 29.341e-18
c1024 n18__ck_buff vss 27.8168e-18
c1025 n20__ck_buff vss 27.6699e-18
c1026 n23__ck_b vss 28.551e-18
c1027 n2__i18__net3 vss 13.785e-18
c1028 n7__i13__net11 vss 103.17e-18
c1029 n7__i13__net12 vss 99.1036e-18
c1030 n2__i13__i19__i4__net2 vss 22.397e-18
c1031 n2__i13__i18__i4__net2 vss 23.5209e-18
c1032 n10__i13__net1 vss 43.7051e-18
c1033 n10__i13__net2 vss 43.6544e-18
c1034 n3__i2__net1 vss 142.801e-18
c1035 n3__i1__net1 vss 146.928e-18
c1036 n3__i0__net1 vss 139.857e-18
c1037 n7__i13__net1 vss 10.089e-18
c1038 n7__i13__net2 vss 9.9191e-18
c1039 n121__i18__net4 vss 21.3111e-18
c1040 n114__i18__net4 vss 15.1524e-18
c1041 n3__i13__i19__net1 vss 50.0268e-18
c1042 n3__i13__i18__net1 vss 51.0698e-18
c1043 n19__shift vss 26.093e-18
c1044 n21__shift vss 26.9882e-18
c1045 n23__shift vss 27.302e-18
c1046 n111__i18__net4 vss 14.8242e-18
c1047 n4__i2__net79 vss 27.2565e-18
c1048 n4__i1__net79 vss 28.5411e-18
c1049 n4__i0__net79 vss 30.968e-18
c1050 n3__i13__net1 vss 25.7831e-18
c1051 n3__i13__net2 vss 23.5841e-18
c1052 n14__shift vss 24.1297e-18
c1053 n16__shift vss 25.5343e-18
c1054 n18__shift vss 23.8564e-18
c1055 n2__i2__net79 vss 28.2511e-18
c1056 n2__i1__net79 vss 30.879e-18
c1057 n2__i0__net79 vss 31.3338e-18
c1058 n104__i18__net4 vss 14.9619e-18
c1059 n3__i13__net11 vss 12.7288e-18
c1060 n3__i13__net12 vss 12.4653e-18
c1061 n3__shift vss 9.11561e-18
c1062 n7__shift vss 9.40393e-18
c1063 n11__shift vss 7.6482e-18
c1064 n101__i18__net4 vss 15.1974e-18
c1065 n96__i18__net4 vss 15.1974e-18
c1066 n89__i18__net4 vss 15.2169e-18
c1067 n12__ck4 vss 47.7132e-18
c1068 n7__i13__a3 vss 101.439e-18
c1069 n7__i13__a1 vss 99.381e-18
c1070 n84__i18__net4 vss 15.2169e-18
c1071 n3__i9__net1 vss 41.9325e-18
c1072 n2__net14 vss 14.5051e-18
c1073 n2__i13__i17__i4__net2 vss 22.3303e-18
c1074 n2__i13__i16__i4__net2 vss 23.4079e-18
c1075 n14__i13__a2 vss 43.5944e-18
c1076 n14__i13__a0 vss 43.5403e-18
c1077 n81__i18__net4 vss 15.2169e-18
c1078 n9__net14 vss 9.34277e-18
c1079 n74__i18__net4 vss 15.2169e-18
c1080 n7__i13__a2 vss 9.9763e-18
c1081 n7__i13__a0 vss 10.0778e-18
c1082 n3__i9__net2 vss 61.3266e-18
c1083 n2__net13 vss 14.8075e-18
c1084 n69__i18__net4 vss 15.1865e-18
c1085 n57__reset vss 6.92224e-18
c1086 n5__i9__i4__net4 vss 19.4364e-18
c1087 n9__net13 vss 8.65283e-18
c1088 n3__i13__i17__net1 vss 50.8335e-18
c1089 n3__i13__i16__net1 vss 50.3137e-18
c1090 n64__i18__net4 vss 15.2169e-18
c1091 n51__reset vss 36.0587e-18
c1092 n60__i18__net4 vss 15.2337e-18
c1093 n3__i13__a2 vss 24.1281e-18
c1094 n3__i13__a0 vss 25.2409e-18
c1095 n28__ck vss 61.1988e-18
c1096 n4__i9__i4__net5 vss 75.0797e-18
c1097 n3__i13__a3 vss 12.1403e-18
c1098 n3__i13__a1 vss 12.1391e-18
c1099 n54__i18__net4 vss 15.2337e-18
c1100 n2__reset_b vss 48.1989e-18
c1101 n49__i18__net4 vss 15.1974e-18
c1102 n46__i18__net4 vss 15.1974e-18
c1103 n41__i18__net4 vss 15.215e-18
c1104 n3__y_out_3 vss 104.467e-18
c1105 n3__y_out_1 vss 101.607e-18
c1106 n3__ck_b vss 25.7823e-18
c1107 n3__ck_buff vss 31.5001e-18
c1108 n38__i18__net4 vss 15.2169e-18
c1109 n2__i13__i15__net2 vss 22.2463e-18
c1110 n2__i13__i13__net2 vss 22.996e-18
c1111 n11__x_out_3 vss 42.4006e-18
c1112 n11__x_out_1 vss 41.8869e-18
c1113 n4__net12 vss 14.568e-18
c1114 n35__i18__net4 vss 15.215e-18
c1115 n4__i9__i4__net1 vss 86.7918e-18
c1116 n8__x_out_3 vss 8.71855e-18
c1117 n8__x_out_1 vss 8.78978e-18
c1118 n32__i18__net4 vss 15.2169e-18
c1119 n29__i18__net4 vss 15.2169e-18
c1120 n26__i18__net4 vss 15.2169e-18
c1121 n23__i18__net4 vss 15.2337e-18
c1122 n3__y_out_2 vss 101.454e-18
c1123 n8__x_out_0 vss 100.032e-18
c1124 n20__i18__net4 vss 15.2033e-18
c1125 n2__i13__i14__net2 vss 22.2594e-18
c1126 n2__i13__i12__net2 vss 23.3336e-18
c1127 n11__x_out_2 vss 38.0062e-18
c1128 n6__y_out_0 vss 38.0168e-18
c1129 n17__i18__net4 vss 15.1974e-18
c1130 n4__net11 vss 13.5206e-18
c1131 n14__i18__net4 vss 15.1974e-18
c1132 n8__x_out_2 vss 9.02754e-18
c1133 n3__y_out_0 vss 8.49964e-18
c1134 n11__i18__net4 vss 15.2169e-18
c1135 n3__i14__x_out_b_1 vss 61.5117e-18
c1136 n3__i14__y_out_b_2 vss 65.0006e-18
c1137 n3__i14__y_out_b_1 vss 66.2444e-18
c1138 n3__i14__x_out_b_0 vss 60.9896e-18
c1139 n8__i18__net4 vss 15.2169e-18
c1140 n8__i14__net7 vss 7.80288e-18
c1141 n8__i14__net11 vss 7.61985e-18
c1142 n5__i18__net4 vss 14.9766e-18
c1143 n5__i14__i11__net4 vss 21.521e-18
c1144 n5__i14__i14__net4 vss 20.7625e-18
c1145 n5__i14__i15__net4 vss 20.6701e-18
c1146 n5__i14__i12__net4 vss 19.5439e-18
c1147 n11__i14__net7 vss 7.79943e-18
c1148 n11__i14__net11 vss 7.18244e-18
c1149 n2__i18__net4 vss 23.187e-18
c1150 n4__i14__i11__net5 vss 75.9042e-18
c1151 n4__i14__i14__net5 vss 79.1708e-18
c1152 n4__i14__i15__net5 vss 76.8183e-18
c1153 n4__i14__i12__net5 vss 73.0119e-18
c1154 n22__i14__net4 vss 46.9241e-18
c1155 n24__i14__net4 vss 46.6306e-18
c1156 n26__i14__net4 vss 46.8345e-18
c1157 n28__i14__net4 vss 45.8401e-18
c1158 n3__i14__net11 vss 117.421e-18
c1159 n32__i14__net4 vss 9.55098e-18
c1160 n3__i14__net7 vss 8.80736e-18
c1161 n35__i14__net4 vss 8.91348e-18
c1162 n57__i14__net10 vss 29.9779e-18
c1163 n49__i14__net9 vss 25.916e-18
c1164 n51__i14__net9 vss 25.916e-18
c1165 n59__i14__net10 vss 30.6737e-18
c1166 n61__i14__net10 vss 30.669e-18
c1167 n53__i14__net9 vss 25.916e-18
c1168 n55__i14__net9 vss 25.916e-18
c1169 n63__i14__net10 vss 30.0956e-18
c1170 n471__i18__net5 vss 20.6999e-18
c1171 n7__i14__i17__net11 vss 30.8956e-18
c1172 n464__i18__net5 vss 15.2214e-18
c1173 n16__i14__i17__net8 vss 30.6251e-18
c1174 n29__reset vss 9.52097e-18
c1175 n5__i14__i17__net11 vss 210.423e-18
c1176 n459__i18__net5 vss 14.8576e-18
c1177 n4__i14__i11__net1 vss 92.8637e-18
c1178 n4__i14__i14__net1 vss 93.7272e-18
c1179 n4__i14__i15__net1 vss 93.7178e-18
c1180 n4__i14__i12__net1 vss 91.4234e-18
c1181 n32__reset vss 6.8751e-18
c1182 n6__i14__i17__net10 vss 52.959e-18
c1183 n29__i14__net3 vss 21.5884e-18
c1184 n31__i14__net3 vss 22.9014e-18
c1185 n33__i14__net3 vss 23.2903e-18
c1186 n35__i14__net3 vss 69.4124e-18
c1187 n454__i18__net5 vss 14.9954e-18
c1188 n451__i18__net5 vss 15.2308e-18
c1189 n6__i14__i17__net9 vss 19.0685e-18
c1190 n3__i14__i17__net9 vss 11.2991e-18
c1191 n444__i18__net5 vss 15.2308e-18
c1192 n12__i14__i17__net8 vss 199.708e-18
c1193 n441__i18__net5 vss 15.2504e-18
c1194 n11__i14__i17__net8 vss 26.2021e-18
c1195 n3__i14__i17__net10 vss 12.6284e-18
c1196 n436__i18__net5 vss 15.2504e-18
c1197 n33__i14__net9 vss 30.1314e-18
c1198 n29__i14__net10 vss 27.7813e-18
c1199 n31__i14__net10 vss 27.7813e-18
c1200 n35__i14__net9 vss 30.5009e-18
c1201 n37__i14__net9 vss 30.5534e-18
c1202 n33__i14__net10 vss 27.7813e-18
c1203 n35__i14__net10 vss 27.7813e-18
c1204 n39__i14__net9 vss 31.367e-18
c1205 n16__i14__i17__net1 vss 57.7029e-18
c1206 n8__i14__i17__net8 vss 60.1874e-18
c1207 n429__i18__net5 vss 15.2504e-18
c1208 n5__i14__i17__i2__net4 vss 19.527e-18
c1209 n5__i14__i17__i3__net4 vss 20.3194e-18
c1210 n3__i14__y_out_b_3 vss 58.8678e-18
c1211 n3__i14__y_out_b_0 vss 59.9779e-18
c1212 n3__i14__x_out_b_2 vss 65.9035e-18
c1213 n3__i14__x_out_b_3 vss 57.9382e-18
c1214 n424__i18__net5 vss 15.2504e-18
c1215 n420__i18__net5 vss 15.2504e-18
c1216 n5__i14__i13__net4 vss 21.2704e-18
c1217 n5__i14__i16__net4 vss 20.8504e-18
c1218 n5__i14__i10__net4 vss 20.8543e-18
c1219 n5__i14__i9__net4 vss 19.8075e-18
c1220 n4__i14__i17__i2__net5 vss 80.5231e-18
c1221 n4__i14__i17__i3__net5 vss 78.234e-18
c1222 n414__i18__net5 vss 15.2504e-18
c1223 n2__i14__i17__net6 vss 44.0272e-18
c1224 n4__i14__i17__net6 vss 47.6594e-18
c1225 n409__i18__net5 vss 15.2671e-18
c1226 n4__i14__i13__net5 vss 80.0285e-18
c1227 n4__i14__i16__net5 vss 78.9246e-18
c1228 n4__i14__i10__net5 vss 82.7728e-18
c1229 n4__i14__i9__net5 vss 76.6136e-18
c1230 n406__i18__net5 vss 15.2671e-18
c1231 n2__i14__net4 vss 45.8126e-18
c1232 n4__i14__net4 vss 45.524e-18
c1233 n6__i14__net4 vss 45.0931e-18
c1234 n8__i14__net4 vss 46.4438e-18
c1235 n399__i18__net5 vss 15.2308e-18
c1236 n6__ck vss 30.5233e-18
c1237 n3__i14__i17__net3 vss 26.8525e-18
c1238 n3__i14__i17__net1 vss 26.6537e-18
c1239 n3__i14__i17__net7 vss 31.2188e-18
c1240 n396__i18__net5 vss 15.2308e-18
c1241 n391__i18__net5 vss 15.2504e-18
c1242 n9__i14__net10 vss 30.0306e-18
c1243 n9__i14__net9 vss 26.0055e-18
c1244 n11__i14__net9 vss 26.0095e-18
c1245 n11__i14__net10 vss 30.6781e-18
c1246 n13__i14__net10 vss 30.673e-18
c1247 n13__i14__net9 vss 26.0122e-18
c1248 n15__i14__net9 vss 26.0082e-18
c1249 n15__i14__net10 vss 31.4909e-18
c1250 n386__i18__net5 vss 15.2504e-18
c1251 n4__i14__i17__i2__net1 vss 91.1051e-18
c1252 n4__i14__i17__i3__net1 vss 89.3343e-18
c1253 n379__i18__net5 vss 15.2504e-18
c1254 n4__reset vss 21.8086e-18
c1255 n6__reset vss 25.4922e-18
c1256 n4__i14__i13__net1 vss 89.6436e-18
c1257 n4__i14__i16__net1 vss 89.9513e-18
c1258 n4__i14__i10__net1 vss 94.5695e-18
c1259 n4__i14__i9__net1 vss 87.4054e-18
c1260 n376__i18__net5 vss 15.2504e-18
c1261 n3__i14__net3 vss 22.8113e-18
c1262 n5__i14__net3 vss 23.2001e-18
c1263 n7__i14__net3 vss 67.6895e-18
c1264 n369__i18__net5 vss 15.2504e-18
c1265 n366__i18__net5 vss 15.2504e-18
c1266 n361__i18__net5 vss 15.2671e-18
c1267 n4__ck vss 25.5669e-18
c1268 n356__i18__net5 vss 15.2671e-18
c1269 n3__i14__net10 vss 29.4931e-18
c1270 n3__i14__net9 vss 32.1228e-18
c1271 n5__i14__net9 vss 32.1677e-18
c1272 n5__i14__net10 vss 29.5632e-18
c1273 n7__i14__net10 vss 29.4931e-18
c1274 n7__i14__net9 vss 31.3955e-18
c1275 n2__ck vss 35.2333e-18
c1276 n2__reset vss 34.0293e-18
c1277 n349__i18__net5 vss 15.2308e-18
c1278 n346__i18__net5 vss 15.2308e-18
c1279 n339__i18__net5 vss 15.2504e-18
c1280 n336__i18__net5 vss 15.2504e-18
c1281 n329__i18__net5 vss 15.2504e-18
c1282 n326__i18__net5 vss 15.2504e-18
c1283 n321__i18__net5 vss 15.2504e-18
c1284 n314__i18__net5 vss 15.2671e-18
c1285 n311__i18__net5 vss 15.2671e-18
c1286 n304__i18__net5 vss 15.2308e-18
c1287 n299__i18__net5 vss 15.2308e-18
c1288 n294__i18__net5 vss 15.2504e-18
c1289 n289__i18__net5 vss 15.2504e-18
c1290 n284__i18__net5 vss 15.2504e-18
c1291 n279__i18__net5 vss 15.2504e-18
c1292 n276__i18__net5 vss 15.2504e-18
c1293 n269__i18__net5 vss 15.2504e-18
c1294 n266__i18__net5 vss 15.2671e-18
c1295 n259__i18__net5 vss 15.2671e-18
c1296 n254__i18__net5 vss 15.2308e-18
c1297 n251__i18__net5 vss 15.2308e-18
c1298 n246__i18__net5 vss 15.2504e-18
c1299 n241__i18__net5 vss 15.2504e-18
c1300 n236__i18__net5 vss 15.2504e-18
c1301 n229__i18__net5 vss 15.2504e-18
c1302 n224__i18__net5 vss 15.2504e-18
c1303 n219__i18__net5 vss 15.2504e-18
c1304 n215__i18__net5 vss 15.2671e-18
c1305 n209__i18__net5 vss 15.2671e-18
c1306 n204__i18__net5 vss 15.2308e-18
c1307 n200__i18__net5 vss 15.2308e-18
c1308 n194__i18__net5 vss 15.2504e-18
c1309 n189__i18__net5 vss 15.2504e-18
c1310 n186__i18__net5 vss 15.2504e-18
c1311 n180__i18__net5 vss 15.2504e-18
c1312 n174__i18__net5 vss 15.2504e-18
c1313 n171__i18__net5 vss 15.2671e-18
c1314 n165__i18__net5 vss 15.2671e-18
c1315 n161__i18__net5 vss 15.2308e-18
c1316 n154__i18__net5 vss 10.6382e-18
c1317 n149__i18__net5 vss 10.6578e-18
c1318 n144__i18__net5 vss 10.6578e-18
c1319 n139__i18__net5 vss 10.6578e-18
c1320 n136__i18__net5 vss 10.6578e-18
c1321 n130__i18__net5 vss 10.6578e-18
c1322 n124__i18__net5 vss 10.7444e-18
c1323 n121__i18__net5 vss 10.6746e-18
c1324 n116__i18__net5 vss 9.81618e-18
c1325 n111__i18__net5 vss 9.72297e-18
c1326 n104__i18__net5 vss 10.6382e-18
c1327 n101__i18__net5 vss 10.6578e-18
c1328 n96__i18__net5 vss 10.6578e-18
c1329 n91__i18__net5 vss 10.6578e-18
c1330 n86__i18__net5 vss 10.6578e-18
c1331 n79__i18__net5 vss 10.6578e-18
c1332 n74__i18__net5 vss 10.6578e-18
c1333 n69__i18__net5 vss 15.2671e-18
c1334 n64__i18__net5 vss 15.2671e-18
c1335 n61__i18__net5 vss 15.2308e-18
c1336 n54__i18__net5 vss 10.6382e-18
c1337 n51__i18__net5 vss 10.6578e-18
c1338 n44__i18__net5 vss 10.6578e-18
c1339 n41__i18__net5 vss 10.6578e-18
c1340 n38__i18__net5 vss 10.6578e-18
c1341 n35__i18__net5 vss 10.6578e-18
c1342 n32__i18__net5 vss 10.6746e-18
c1343 n29__i18__net5 vss 10.6746e-18
c1344 n26__i18__net5 vss 10.6382e-18
c1345 n23__i18__net5 vss 10.6382e-18
c1346 n20__i18__net5 vss 10.6578e-18
c1347 n17__i18__net5 vss 10.6578e-18
c1348 n14__i18__net5 vss 10.6578e-18
c1349 n11__i18__net5 vss 10.6578e-18
c1350 n8__i18__net5 vss 10.6578e-18
c1351 n5__i18__net5 vss 10.4174e-18
c1352 n2__i18__net5 vss 19.3564e-18
c1353 n1021__vddio vss 125.658e-18
c1354 n30__vdd vss 1.00275e-15
c1355 n439__vddio vss 825.048e-18
c1356 n19__vdd vss 1.76839e-15
c1357 n458__r_out vss 650.746e-18
c1358 n1010__vddio vss 151.251e-18
c1359 n1011__vddio vss 706.319e-18
c1360 n1012__vddio vss 380.796e-18
c1361 n1013__vddio vss 191.39e-18
c1362 n1014__vddio vss 121.429e-18
c1363 n1015__vddio vss 18.9027e-18
c1364 n1016__vddio vss 9.13519e-18
c1365 n29__vdd vss 221.538e-18
c1366 n435__vddio vss 49.0147e-18
c1367 n436__vddio vss 72.0154e-18
c1368 n437__vddio vss 48.4182e-18
c1369 n438__vddio vss 4.55949e-18
c1370 n14__vdd vss 54.8206e-18
c1371 n15__vdd vss 93.4839e-18
c1372 n18__vdd vss 153.194e-18
c1373 n459__r_out vss 2.58979e-18
c1374 n1003__vddio vss 3.68024e-18
c1375 n1004__vddio vss 2.17024e-18
c1376 n1005__vddio vss 2.28797e-18
c1377 n1006__vddio vss 2.28797e-18
c1378 n1007__vddio vss 2.28797e-18
c1379 n1008__vddio vss 2.16725e-18
c1380 n1009__vddio vss 2.28797e-18
c1381 n427__vdd vss 140.752e-18
c1382 n428__vdd vss 152.724e-18
c1383 n28__vdd vss 2.17426e-18
c1384 n13__vdd vss 726.635e-21
c1385 n17__vdd vss 93.676e-21
c1386 n996__vddio vss 17.4525e-18
c1387 n998__vddio vss 2.16725e-18
c1388 n999__vddio vss 2.16725e-18
c1389 n1000__vddio vss 2.16725e-18
c1390 n1002__vddio vss 2.16725e-18
c1391 n425__vdd vss 31.3464e-18
c1392 n430__r_out vss 4.20247e-18
c1393 n990__vddio vss 28.5541e-18
c1394 n424__vdd vss 20.1501e-18
c1395 n26__vdd vss 6.14521e-18
c1396 n66__reset vss 169.613e-18
c1397 n37__ck vss 44.8369e-18
c1398 n59__reset vss 196.382e-18
c1399 n33__ck vss 397.445e-18
c1400 n50__reset vss 577.702e-18
c1401 n10__vdd vss 46.0333e-18
c1402 n11__vdd vss 29.482e-18
c1403 n12__vdd vss 29.482e-18
c1404 n20__ck vss 348.709e-18
c1405 n431__r_out vss 33.5766e-18
c1406 n16__r0_buff vss 1.00259e-15
c1407 n17__r2_buff vss 953.796e-18
c1408 n16__r1_buff vss 1.55768e-15
c1409 n976__vddio vss 27.6511e-18
c1410 n977__vddio vss 24.0672e-18
c1411 n17__serial_out_b_high vss 125.525e-18
c1412 n31__serial_out vss 170.614e-18
c1413 n32__serial_out vss 203.218e-18
c1414 n421__vdd vss 39.3567e-18
c1415 n422__vdd vss 39.9842e-18
c1416 n30__serial_out vss 142.798e-18
c1417 n29__serial_out vss 43.0611e-18
c1418 n17__net4 vss 223.632e-18
c1419 n15__net3 vss 295.989e-18
c1420 n16__serial_out_b_high vss 115.542e-18
c1421 n205__i18__net4 vss 26.2074e-18
c1422 n206__i18__net4 vss 56.7497e-18
c1423 n194__i18__net4 vss 38.3947e-18
c1424 n195__i18__net4 vss 49.7241e-18
c1425 n174__i18__net4 vss 37.9201e-18
c1426 n177__i18__net4 vss 48.6676e-18
c1427 n172__i18__net4 vss 38.265e-18
c1428 n173__i18__net4 vss 48.8309e-18
c1429 n161__i18__net4 vss 85.057e-18
c1430 n162__i18__net4 vss 130.093e-18
c1431 n21__reset_b vss 642.323e-18
c1432 n37__ck_buff vss 229.708e-18
c1433 n28__reset_buff vss 352.113e-18
c1434 n31__ck_b vss 783.056e-18
c1435 n695__i18__net5 vss 37.1329e-18
c1436 n696__i18__net5 vss 24.3351e-18
c1437 n6__net4 vss 126.379e-18
c1438 n7__net4 vss 333.75e-18
c1439 n25__vdd vss 18.7339e-18
c1440 n7__r0_buff vss 119.891e-18
c1441 n7__r1_buff vss 178.069e-18
c1442 n7__r2_buff vss 168.866e-18
c1443 n675__i18__net5 vss 38.7274e-18
c1444 n676__i18__net5 vss 51.0059e-18
c1445 n3__net4 vss 112.96e-18
c1446 n3__net3 vss 373.162e-18
c1447 n669__i18__net5 vss 38.7847e-18
c1448 n670__i18__net5 vss 49.7059e-18
c1449 n2__r2_buff vss 1.26334e-15
c1450 n19__reset_buff vss 246.155e-18
c1451 n2__r1_buff vss 1.7692e-15
c1452 n656__i18__net5 vss 41.1907e-18
c1453 n657__i18__net5 vss 39.1646e-18
c1454 n2__r0_buff vss 1.46463e-15
c1455 n632__i18__net5 vss 38.7655e-18
c1456 n635__i18__net5 vss 50.0509e-18
c1457 n23__ck_buff vss 432.868e-18
c1458 n630__i18__net5 vss 41.2648e-18
c1459 n631__i18__net5 vss 40.4956e-18
c1460 n62__reset vss 28.2037e-18
c1461 n617__i18__net5 vss 39.0838e-18
c1462 n618__i18__net5 vss 52.1474e-18
c1463 n36__ck vss 47.8216e-18
c1464 n21__i13__a2 vss 86.8148e-18
c1465 n22__i13__a0 vss 89.3072e-18
c1466 n597__i18__net5 vss 38.8724e-18
c1467 n598__i18__net5 vss 48.7197e-18
c1468 n591__i18__net5 vss 39.2547e-18
c1469 n592__i18__net5 vss 51.717e-18
c1470 n20__x_out_1 vss 389.175e-18
c1471 n21__x_out_1 vss 188.95e-18
c1472 n15__y_out_1 vss 385.412e-18
c1473 n16__y_out_1 vss 185.18e-18
c1474 n32__ck vss 53.1893e-18
c1475 n10__y_out_3 vss 487.395e-18
c1476 n11__y_out_3 vss 351.365e-18
c1477 n10__y_out_1 vss 50.6983e-18
c1478 n578__i18__net5 vss 39.1779e-18
c1479 n579__i18__net5 vss 38.4853e-18
c1480 n8__reset_buff vss 55.4192e-18
c1481 n9__reset_buff vss 164.401e-18
c1482 n14__x_out_3 vss 534.164e-18
c1483 n15__x_out_1 vss 65.8745e-18
c1484 n7__reset_buff vss 50.9946e-18
c1485 n19__i13__a2 vss 188.342e-18
c1486 n20__i13__a0 vss 143.164e-18
c1487 n558__i18__net5 vss 39.7379e-18
c1488 n559__i18__net5 vss 54.5937e-18
c1489 n5__reset_b vss 605.266e-18
c1490 n3__reset_b vss 39.5561e-18
c1491 n8__ck_buff vss 325.369e-18
c1492 n15__ck_b vss 731.151e-18
c1493 n552__i18__net5 vss 38.6919e-18
c1494 n553__i18__net5 vss 52.1493e-18
c1495 n15__y_out_2 vss 231.546e-18
c1496 n16__y_out_2 vss 107.364e-18
c1497 n19__x_out_2 vss 330.574e-18
c1498 n20__x_out_2 vss 144.979e-18
c1499 n539__i18__net5 vss 38.5233e-18
c1500 n540__i18__net5 vss 50.8889e-18
c1501 n10__y_out_2 vss 61.7505e-18
c1502 n13__x_out_0 vss 215.843e-18
c1503 n15__x_out_2 vss 91.6443e-18
c1504 n13__y_out_0 vss 102e-18
c1505 n109__i14__net10 vss 676.563e-18
c1506 n110__i14__net10 vss 704.224e-18
c1507 n111__i14__net10 vss 713.954e-18
c1508 n112__i14__net10 vss 617.506e-18
c1509 n526__i18__net5 vss 39.0892e-18
c1510 n527__i18__net5 vss 52.0245e-18
c1511 n5__y_out_3 vss 251.293e-18
c1512 n6__y_out_2 vss 132.966e-18
c1513 n5__y_out_1 vss 317.473e-18
c1514 n8__y_out_0 vss 81.0292e-18
c1515 n39__i14__net7 vss 66.3355e-18
c1516 n38__i14__net11 vss 24.3572e-18
c1517 n513__i18__net5 vss 77.081e-18
c1518 n514__i18__net5 vss 133.586e-18
c1519 n36__i14__net7 vss 151.71e-18
c1520 n35__i14__net11 vss 64.4059e-18
c1521 n12__x_out_3 vss 408.499e-18
c1522 n13__x_out_3 vss 469.779e-18
c1523 n12__x_out_2 vss 469.612e-18
c1524 n13__x_out_2 vss 222.472e-18
c1525 n12__x_out_1 vss 465.061e-18
c1526 n13__x_out_1 vss 469.775e-18
c1527 n10__x_out_0 vss 473.346e-18
c1528 n11__x_out_0 vss 197.153e-18
c1529 n82__i14__net9 vss 592.318e-18
c1530 n83__i14__net9 vss 537.959e-18
c1531 n84__i14__net9 vss 533.534e-18
c1532 n85__i14__net9 vss 499.1e-18
c1533 n64__i14__net3 vss 360.759e-18
c1534 n65__i14__net3 vss 372.261e-18
c1535 n66__i14__net3 vss 371.386e-18
c1536 n67__i14__net3 vss 343.545e-18
c1537 n31__i14__net7 vss 154.12e-18
c1538 n29__i14__net11 vss 149.274e-18
c1539 n68__i14__net4 vss 509.326e-18
c1540 n654__r_out vss 24.6989e-18
c1541 n655__r_out vss 37.554e-18
c1542 n641__r_out vss 41.906e-18
c1543 n642__r_out vss 61.0163e-18
c1544 n53__i14__net3 vss 1.03597e-15
c1545 n54__i14__net3 vss 1.03547e-15
c1546 n55__i14__net3 vss 1.05019e-15
c1547 n56__i14__net3 vss 1.05412e-15
c1548 n47__reset vss 383.511e-18
c1549 n89__i14__net10 vss 1.11471e-15
c1550 n90__i14__net10 vss 1.1143e-15
c1551 n91__i14__net10 vss 1.13536e-15
c1552 n92__i14__net10 vss 1.13495e-15
c1553 n628__r_out vss 39.2816e-18
c1554 n629__r_out vss 44.2117e-18
c1555 n69__i14__net9 vss 1.11054e-15
c1556 n70__i14__net9 vss 1.10898e-15
c1557 n71__i14__net9 vss 1.11395e-15
c1558 n72__i14__net9 vss 1.10888e-15
c1559 n615__r_out vss 40.1639e-18
c1560 n616__r_out vss 45.361e-18
c1561 n16__i14__i17__net7 vss 142.694e-18
c1562 n4__y3 vss 478.74e-18
c1563 n5__y2 vss 517.674e-18
c1564 n4__y1 vss 517.556e-18
c1565 n5__y0 vss 467.56e-18
c1566 n25__i14__i17__net1 vss 102.388e-18
c1567 n5__x_out_3 vss 427.747e-18
c1568 n5__x_out_2 vss 427.764e-18
c1569 n5__x_out_1 vss 427.746e-18
c1570 n5__x_out_0 vss 427.766e-18
c1571 n602__r_out vss 39.7496e-18
c1572 n603__r_out vss 60.1272e-18
c1573 n21__i14__i17__net1 vss 88.4489e-18
c1574 n22__i14__i17__net1 vss 250.771e-18
c1575 n587__r_out vss 39.9609e-18
c1576 n590__r_out vss 41.5962e-18
c1577 n13__i14__i17__net7 vss 98.0436e-18
c1578 n14__i14__i17__net7 vss 257.934e-18
c1579 n576__r_out vss 40.2113e-18
c1580 n577__r_out vss 60.7208e-18
c1581 n9__i14__net4 vss 689.122e-18
c1582 n12__i14__net4 vss 684.648e-18
c1583 n13__i14__net4 vss 698.356e-18
c1584 n16__i14__net4 vss 705.544e-18
c1585 n7__vdd vss 32.939e-18
c1586 n8__vdd vss 36.5166e-18
c1587 n9__vdd vss 36.3972e-18
c1588 n563__r_out vss 39.8802e-18
c1589 n564__r_out vss 46.4761e-18
c1590 n550__r_out vss 38.7041e-18
c1591 n551__r_out vss 45.3626e-18
c1592 n25__reset vss 279.946e-18
c1593 n537__r_out vss 40.1158e-18
c1594 n538__r_out vss 57.7707e-18
c1595 n19__ck vss 13.0755e-18
c1596 n17__i14__net3 vss 665.731e-18
c1597 n18__i14__net3 vss 667.556e-18
c1598 n19__i14__net3 vss 686.887e-18
c1599 n20__i14__net3 vss 684.311e-18
c1600 n524__r_out vss 41.7212e-18
c1601 n525__r_out vss 41.9309e-18
c1602 n45__i14__net10 vss 243.687e-18
c1603 n46__i14__net10 vss 243.351e-18
c1604 n47__i14__net10 vss 260.953e-18
c1605 n48__i14__net10 vss 260.28e-18
c1606 n9__i14__i17__net7 vss 217.858e-18
c1607 n29__i14__net9 vss 520.883e-18
c1608 n30__i14__net9 vss 520.876e-18
c1609 n31__i14__net9 vss 546.481e-18
c1610 n32__i14__net9 vss 539.491e-18
c1611 n12__i14__i17__net1 vss 285.435e-18
c1612 n504__r_out vss 39.888e-18
c1613 n505__r_out vss 61.255e-18
c1614 n13__reset vss 485.621e-18
c1615 n5__x3 vss 7.50814e-18
c1616 n5__x2 vss 7.3997e-18
c1617 n5__x1 vss 25.518e-18
c1618 n5__x0 vss 25.4928e-18
c1619 n491__r_out vss 39.6848e-18
c1620 n492__r_out vss 45.5273e-18
c1621 n485__r_out vss 40.1667e-18
c1622 n486__r_out vss 45.361e-18
c1623 n472__r_out vss 40.3889e-18
c1624 n473__r_out vss 63.1175e-18
c1625 n456__r_out vss 40.1311e-18
c1626 n457__r_out vss 41.4818e-18
c1627 n436__r_out vss 39.4325e-18
c1628 n437__r_out vss 58.86e-18
c1629 n428__r_out vss 39.8535e-18
c1630 n429__r_out vss 45.4915e-18
c1631 n415__r_out vss 40.4588e-18
c1632 n416__r_out vss 45.2553e-18
c1633 n402__r_out vss 39.6828e-18
c1634 n403__r_out vss 61.1481e-18
c1635 n389__r_out vss 39.8022e-18
c1636 n390__r_out vss 41.3944e-18
c1637 n369__r_out vss 40.2306e-18
c1638 n370__r_out vss 63.0658e-18
c1639 n363__r_out vss 39.7519e-18
c1640 n364__r_out vss 44.0698e-18
c1641 n350__r_out vss 39.5531e-18
c1642 n351__r_out vss 45.2814e-18
c1643 n330__r_out vss 40.1915e-18
c1644 n331__r_out vss 60.0918e-18
c1645 n317__r_out vss 40.4567e-18
c1646 n318__r_out vss 41.7094e-18
c1647 n304__r_out vss 39.9072e-18
c1648 n305__r_out vss 61.4958e-18
c1649 n291__r_out vss 39.7042e-18
c1650 n292__r_out vss 45.5571e-18
c1651 n285__r_out vss 40.1576e-18
c1652 n286__r_out vss 45.0999e-18
c1653 n265__r_out vss 40.2284e-18
c1654 n266__r_out vss 63.0359e-18
c1655 n252__r_out vss 39.9536e-18
c1656 n253__r_out vss 41.4017e-18
c1657 n239__r_out vss 39.4325e-18
c1658 n240__r_out vss 53.1691e-18
c1659 n226__r_out vss 39.8535e-18
c1660 n227__r_out vss 39.3328e-18
c1661 n220__r_out vss 40.4588e-18
c1662 n221__r_out vss 37.9373e-18
c1663 n200__r_out vss 39.9193e-18
c1664 n201__r_out vss 51.1193e-18
c1665 n194__r_out vss 22.2816e-18
c1666 n195__r_out vss 20.5586e-18
c1667 n174__r_out vss 21.7807e-18
c1668 n175__r_out vss 38.8614e-18
c1669 n168__r_out vss 39.8409e-18
c1670 n169__r_out vss 38.6501e-18
c1671 n155__r_out vss 39.6704e-18
c1672 n156__r_out vss 37.3337e-18
c1673 n142__r_out vss 40.1069e-18
c1674 n143__r_out vss 50.6079e-18
c1675 n122__r_out vss 40.4567e-18
c1676 n123__r_out vss 43.3076e-18
c1677 n109__r_out vss 39.9072e-18
c1678 n110__r_out vss 62.3927e-18
c1679 n96__r_out vss 39.684e-18
c1680 n97__r_out vss 45.9103e-18
c1681 n90__r_out vss 40.1374e-18
c1682 n91__r_out vss 48.2468e-18
c1683 n70__r_out vss 40.0506e-18
c1684 n71__r_out vss 59.6742e-18
c1685 n64__r_out vss 39.8702e-18
c1686 n65__r_out vss 43.7618e-18
c1687 n44__r_out vss 39.4378e-18
c1688 n45__r_out vss 58.0815e-18
c1689 n38__r_out vss 39.777e-18
c1690 n39__r_out vss 47.3378e-18
c1691 n25__r_out vss 40.4671e-18
c1692 n26__r_out vss 47.8701e-18
c1693 n5__r_out vss 160.034e-18
c1694 n6__r_out vss 138.889e-18
c1695 n970__vddio vss 20.2114e-18
c1696 n971__vddio vss 10.1412e-18
c1697 n972__vddio vss 10.1412e-18
c1698 n973__vddio vss 7.81891e-18
c1699 n974__vddio vss 3.69276e-18
c1700 n15__serial_out_b_high vss 22.0994e-18
c1701 n968__vddio vss 100.927e-18
c1702 n10__r2 vss 490.074e-18
c1703 n15__r0 vss 466.839e-18
c1704 n15__r1 vss 268.078e-18
c1705 n26__serial_out vss 286.282e-18
c1706 n967__vddio vss 89.8493e-18
c1707 n25__serial_out vss 50.1907e-18
c1708 n16__net4 vss 81.0511e-18
c1709 n14__net3 vss 50.2046e-18
c1710 n14__serial_out_b_high vss 115.125e-18
c1711 n50__i18__net3 vss 5.67233e-18
c1712 n203__i18__net4 vss 12.1981e-18
c1713 n204__i18__net4 vss 8.77955e-18
c1714 n48__i18__net3 vss 9.41857e-18
c1715 n966__vddio vss 5.30089e-18
c1716 n47__i18__net3 vss 9.41857e-18
c1717 n192__i18__net4 vss 9.58205e-18
c1718 n193__i18__net4 vss 7.20114e-18
c1719 n44__i18__net3 vss 9.20133e-18
c1720 n4__r2 vss 459.607e-18
c1721 n42__i18__net3 vss 9.20133e-18
c1722 n11__i13__net23 vss 477.371e-18
c1723 n10__i13__net23 vss 180.875e-18
c1724 n175__i18__net4 vss 3.15399e-18
c1725 n176__i18__net4 vss 6.84019e-18
c1726 n40__i18__net3 vss 9.30995e-18
c1727 n38__i18__net3 vss 9.30995e-18
c1728 n170__i18__net4 vss 2.07787e-18
c1729 n171__i18__net4 vss 7.07967e-18
c1730 n37__i18__net3 vss 9.30995e-18
c1731 n10__i13__net17 vss 261.96e-18
c1732 n11__i13__net17 vss 148.522e-18
c1733 n13__i13__net7 vss 224.521e-18
c1734 n15__i13__net7 vss 218.123e-18
c1735 n34__i18__net3 vss 9.88756e-18
c1736 n21__i13__net18 vss 110.593e-18
c1737 n19__i13__net18 vss 105.25e-18
c1738 n159__i18__net4 vss 11.5669e-18
c1739 n9__r0 vss 519.508e-18
c1740 n32__i18__net3 vss 12.1121e-18
c1741 n22__reset_b vss 513.869e-18
c1742 n23__reset_b vss 602.032e-18
c1743 n24__reset_b vss 531.943e-18
c1744 n34__ck_buff vss 365.191e-18
c1745 n36__ck_buff vss 311.579e-18
c1746 n35__ck_buff vss 179.494e-18
c1747 n26__reset_buff vss 494.022e-18
c1748 n27__reset_buff vss 495.899e-18
c1749 n29__reset_buff vss 517.216e-18
c1750 n633__vddio vss 283.106e-18
c1751 n634__vddio vss 80.1519e-18
c1752 n635__vddio vss 10.4155e-18
c1753 n626__vddio vss 11.431e-18
c1754 n150__i18__net4 vss 26.0782e-18
c1755 n32__ck_b vss 282.464e-18
c1756 n33__ck_b vss 390.093e-18
c1757 n34__ck_b vss 261.683e-18
c1758 n694__i18__net5 vss 26.6119e-18
c1759 n148__i18__net4 vss 8.66091e-18
c1760 n6__r0_buff vss 99.0348e-18
c1761 n6__r1_buff vss 97.8095e-18
c1762 n6__r2_buff vss 84.7149e-18
c1763 n530__vddio vss 63.362e-18
c1764 n531__vddio vss 39.0283e-18
c1765 n534__vddio vss 21.8548e-18
c1766 n146__i18__net4 vss 9.41857e-18
c1767 n671__i18__net5 vss 9.58205e-18
c1768 n674__i18__net5 vss 7.2635e-18
c1769 n2__net3 vss 115.729e-18
c1770 n144__i18__net4 vss 9.41857e-18
c1771 n524__vddio vss 62.7713e-18
c1772 n525__vddio vss 36.8858e-18
c1773 n528__vddio vss 20.3568e-18
c1774 n142__i18__net4 vss 9.20133e-18
c1775 n13__i13__net11 vss 159.126e-18
c1776 n14__i13__net11 vss 86.2938e-18
c1777 n19__i13__net2 vss 96.6354e-18
c1778 n20__i13__net2 vss 77.0752e-18
c1779 n667__i18__net5 vss 8.90714e-18
c1780 n15__i13__net1 vss 211.937e-18
c1781 n17__i13__net12 vss 154.718e-18
c1782 n18__i13__net12 vss 175.221e-18
c1783 n140__i18__net4 vss 9.20133e-18
c1784 n16__i13__net1 vss 280.504e-18
c1785 n518__vddio vss 56.6799e-18
c1786 n519__vddio vss 34.463e-18
c1787 n522__vddio vss 19.0098e-18
c1788 n138__i18__net4 vss 9.30995e-18
c1789 n16__reset_buff vss 138.461e-18
c1790 n17__ck4 vss 258.624e-18
c1791 n655__i18__net5 vss 17.6735e-18
c1792 n136__i18__net4 vss 9.30995e-18
c1793 n512__vddio vss 57.1345e-18
c1794 n513__vddio vss 34.463e-18
c1795 n516__vddio vss 19.0098e-18
c1796 n134__i18__net4 vss 9.30995e-18
c1797 n633__i18__net5 vss 3.50388e-18
c1798 n634__i18__net5 vss 6.88309e-18
c1799 n132__i18__net4 vss 9.30995e-18
c1800 n22__ck_buff vss 37.4361e-18
c1801 n505__vddio vss 63.4345e-18
c1802 n508__vddio vss 28.2259e-18
c1803 n509__vddio vss 24.0596e-18
c1804 n130__i18__net4 vss 9.30995e-18
c1805 n64__reset vss 9.60176e-18
c1806 n628__i18__net5 vss 5.91466e-18
c1807 n629__i18__net5 vss 10.6675e-18
c1808 n128__i18__net4 vss 9.30995e-18
c1809 n61__reset vss 8.82839e-18
c1810 n499__vddio vss 55.3117e-18
c1811 n502__vddio vss 34.3673e-18
c1812 n503__vddio vss 24.3758e-18
c1813 n126__i18__net4 vss 9.41857e-18
c1814 n615__i18__net5 vss 3.82761e-18
c1815 n616__i18__net5 vss 7.16768e-18
c1816 n124__i18__net4 vss 9.41857e-18
c1817 n494__vddio vss 63.3235e-18
c1818 n495__vddio vss 37.8824e-18
c1819 n498__vddio vss 20.8763e-18
c1820 n22__i13__a2 vss 66.2028e-18
c1821 n18__i13__a3 vss 45.4487e-18
c1822 n17__i13__a3 vss 40.0221e-18
c1823 n17__i13__a1 vss 39.9115e-18
c1824 n18__i13__a1 vss 45.3731e-18
c1825 n21__i13__a0 vss 66.3228e-18
c1826 n630__vddio vss 14.758e-18
c1827 n118__i18__net4 vss 9.20133e-18
c1828 n594__i18__net5 vss 8.89584e-18
c1829 n117__i18__net4 vss 9.20133e-18
c1830 n488__vddio vss 60.2778e-18
c1831 n489__vddio vss 37.2891e-18
c1832 n492__vddio vss 19.9554e-18
c1833 n109__i18__net4 vss 9.30995e-18
c1834 n589__i18__net5 vss 2.05364e-18
c1835 n590__i18__net5 vss 7.0688e-18
c1836 n107__i18__net4 vss 9.30995e-18
c1837 n482__vddio vss 58.0037e-18
c1838 n483__vddio vss 34.7065e-18
c1839 n486__vddio vss 18.5938e-18
c1840 n99__i18__net4 vss 9.30995e-18
c1841 n12__y_out_3 vss 75.795e-18
c1842 n11__y_out_1 vss 78.3716e-18
c1843 n576__i18__net5 vss 3.55191e-18
c1844 n577__i18__net5 vss 20.0475e-18
c1845 n93__i18__net4 vss 9.30995e-18
c1846 n15__x_out_3 vss 331.43e-18
c1847 n14__x_out_1 vss 94.0601e-18
c1848 n476__vddio vss 51.0539e-18
c1849 n477__vddio vss 31.5424e-18
c1850 n480__vddio vss 17.0509e-18
c1851 n6__reset_buff vss 538.673e-18
c1852 n20__i13__a2 vss 58.643e-18
c1853 n19__i13__a0 vss 62.8451e-18
c1854 n92__i18__net4 vss 9.30995e-18
c1855 n555__i18__net5 vss 7.99099e-18
c1856 n6__reset_b vss 422.906e-18
c1857 n4__reset_b vss 72.3705e-18
c1858 n87__i18__net4 vss 9.30995e-18
c1859 n9__ck_buff vss 194.949e-18
c1860 n470__vddio vss 55.4132e-18
c1861 n471__vddio vss 33.1388e-18
c1862 n474__vddio vss 18.2006e-18
c1863 n632__vddio vss 15.3777e-18
c1864 n79__i18__net4 vss 9.41857e-18
c1865 n550__i18__net5 vss 9.55425e-18
c1866 n551__i18__net5 vss 7.16425e-18
c1867 n77__i18__net4 vss 9.41857e-18
c1868 n464__vddio vss 63.0201e-18
c1869 n465__vddio vss 37.9207e-18
c1870 n468__vddio vss 20.9631e-18
c1871 n72__i18__net4 vss 9.20133e-18
c1872 n12__ck_b vss 62.2297e-18
c1873 n537__i18__net5 vss 3.16692e-18
c1874 n538__i18__net5 vss 6.81202e-18
c1875 n9__ck4 vss 450.082e-18
c1876 n11__y_out_2 vss 104.265e-18
c1877 n12__x_out_0 vss 95.5596e-18
c1878 n67__i18__net4 vss 9.20133e-18
c1879 n14__ck_b vss 99.1147e-18
c1880 n14__x_out_2 vss 59.9504e-18
c1881 n12__y_out_0 vss 41.1034e-18
c1882 n457__vddio vss 71.0622e-18
c1883 n460__vddio vss 31.5509e-18
c1884 n461__vddio vss 27.3894e-18
c1885 n5__ck4 vss 146.812e-18
c1886 n62__i18__net4 vss 9.30995e-18
c1887 n106__i14__net10 vss 53.0399e-18
c1888 n524__i18__net5 vss 2.05364e-18
c1889 n525__i18__net5 vss 7.05163e-18
c1890 n6__y_out_3 vss 67.9175e-18
c1891 n5__y_out_2 vss 64.7517e-18
c1892 n6__y_out_1 vss 21.5838e-18
c1893 n7__y_out_0 vss 20.9354e-18
c1894 n57__i18__net4 vss 9.30995e-18
c1895 n451__vddio vss 66.0482e-18
c1896 n454__vddio vss 29.3098e-18
c1897 n455__vddio vss 24.9532e-18
c1898 n52__i18__net4 vss 9.30995e-18
c1899 n503__i18__net5 vss 11.885e-18
c1900 n35__i14__net7 vss 56.7188e-18
c1901 n44__i18__net4 vss 16.7659e-18
c1902 n430__vddio vss 45.5176e-18
c1903 n431__vddio vss 18.421e-18
c1904 n434__vddio vss 9.93546e-18
c1905 n81__i14__net9 vss 121.956e-18
c1906 n413__vddio vss 17.5961e-18
c1907 n414__vddio vss 3.98298e-18
c1908 n415__vddio vss 3.97648e-18
c1909 n416__vddio vss 2.49451e-18
c1910 n63__i14__net3 vss 84.96e-18
c1911 n30__i14__net11 vss 261.615e-18
c1912 n58__i14__net4 vss 135.874e-18
c1913 n61__i14__net4 vss 188.44e-18
c1914 n62__i14__net4 vss 1.02006e-15
c1915 n64__i14__net4 vss 951.422e-18
c1916 n66__i14__net4 vss 951.325e-18
c1917 n69__i14__net4 vss 492.658e-18
c1918 n401__vddio vss 27.7946e-18
c1919 n404__vddio vss 13.5414e-18
c1920 n405__vddio vss 12.1432e-18
c1921 n408__vddio vss 7.95952e-18
c1922 n500__i18__net5 vss 40.635e-18
c1923 n652__r_out vss 12.1798e-18
c1924 n653__r_out vss 8.50823e-18
c1925 n498__i18__net5 vss 8.99592e-18
c1926 n393__vddio vss 65.6688e-18
c1927 n396__vddio vss 28.7833e-18
c1928 n397__vddio vss 26.0543e-18
c1929 n400__vddio vss 17.344e-18
c1930 n496__i18__net5 vss 10.6368e-18
c1931 n639__r_out vss 3.49208e-18
c1932 n640__r_out vss 6.88871e-18
c1933 n49__i14__net3 vss 20.0035e-18
c1934 n50__i14__net3 vss 517.064e-18
c1935 n51__i14__net3 vss 502.88e-18
c1936 n52__i14__net3 vss 501.373e-18
c1937 n494__i18__net5 vss 9.41857e-18
c1938 n386__vddio vss 62.6458e-18
c1939 n387__vddio vss 37.4089e-18
c1940 n390__vddio vss 22.2861e-18
c1941 n391__vddio vss 13.0382e-18
c1942 n46__reset vss 99.133e-18
c1943 n492__i18__net5 vss 9.20133e-18
c1944 n626__r_out vss 3.16647e-18
c1945 n627__r_out vss 6.5295e-18
c1946 n12__i14__i17__net9 vss 107.317e-18
c1947 n13__i14__i17__net9 vss 120.159e-18
c1948 n61__i14__net9 vss 265.488e-18
c1949 n65__i14__net9 vss 266.183e-18
c1950 n490__i18__net5 vss 9.20133e-18
c1951 n377__vddio vss 71.5393e-18
c1952 n380__vddio vss 31.575e-18
c1953 n381__vddio vss 29.2381e-18
c1954 n384__vddio vss 20.0031e-18
c1955 n488__i18__net5 vss 9.30995e-18
c1956 n8__i14__i17__net10 vss 145.502e-18
c1957 n10__i14__i17__net10 vss 206.196e-18
c1958 n613__r_out vss 2.08912e-18
c1959 n486__i18__net5 vss 9.30995e-18
c1960 n15__i14__i17__net7 vss 103.821e-18
c1961 n8__i14__i17__net11 vss 100.606e-18
c1962 n9__i14__i17__net11 vss 108.334e-18
c1963 n369__vddio vss 67.9408e-18
c1964 n372__vddio vss 30.1552e-18
c1965 n373__vddio vss 27.4767e-18
c1966 n376__vddio vss 18.5992e-18
c1967 n5__y3 vss 49.2897e-18
c1968 n4__y2 vss 49.2197e-18
c1969 n5__y1 vss 152.331e-18
c1970 n4__y0 vss 152.327e-18
c1971 n484__i18__net5 vss 9.30995e-18
c1972 n23__i14__i17__net1 vss 335.499e-18
c1973 n24__i14__i17__net1 vss 44.3681e-18
c1974 n18__i14__i17__net8 vss 76.6442e-18
c1975 n17__i14__i17__net8 vss 361.898e-18
c1976 n4__x_out_3 vss 54.2425e-18
c1977 n4__x_out_2 vss 54.4771e-18
c1978 n4__x_out_1 vss 87.7843e-18
c1979 n4__x_out_0 vss 84.8063e-18
c1980 n600__r_out vss 3.51592e-18
c1981 n601__r_out vss 6.58267e-18
c1982 n482__i18__net5 vss 9.30995e-18
c1983 n361__vddio vss 68.4371e-18
c1984 n364__vddio vss 30.1552e-18
c1985 n365__vddio vss 27.4767e-18
c1986 n368__vddio vss 18.5774e-18
c1987 n480__i18__net5 vss 9.30995e-18
c1988 n588__r_out vss 8.08148e-18
c1989 n478__i18__net5 vss 9.30995e-18
c1990 n353__vddio vss 66.2711e-18
c1991 n356__vddio vss 29.3337e-18
c1992 n357__vddio vss 26.7873e-18
c1993 n360__vddio vss 17.9945e-18
c1994 n476__i18__net5 vss 9.41857e-18
c1995 n574__r_out vss 3.48342e-18
c1996 n575__r_out vss 6.87191e-18
c1997 n474__i18__net5 vss 9.41857e-18
c1998 n346__vddio vss 59.8396e-18
c1999 n347__vddio vss 35.8758e-18
c2000 n350__vddio vss 21.9749e-18
c2001 n351__vddio vss 13.2577e-18
c2002 n10__i14__net4 vss 729.021e-18
c2003 n11__i14__net4 vss 527.448e-18
c2004 n14__i14__net4 vss 546.083e-18
c2005 n15__i14__net4 vss 553.924e-18
c2006 n469__i18__net5 vss 9.20133e-18
c2007 n2__vdd vss 26.7413e-18
c2008 n3__vdd vss 23.962e-18
c2009 n6__vdd vss 23.4207e-18
c2010 n561__r_out vss 3.17923e-18
c2011 n562__r_out vss 6.7225e-18
c2012 n466__i18__net5 vss 9.20133e-18
c2013 n337__vddio vss 72.4332e-18
c2014 n340__vddio vss 32.4552e-18
c2015 n341__vddio vss 30.2336e-18
c2016 n344__vddio vss 21.0052e-18
c2017 n462__i18__net5 vss 9.30995e-18
c2018 n548__r_out vss 2.06465e-18
c2019 n549__r_out vss 6.82799e-18
c2020 n457__i18__net5 vss 9.30995e-18
c2021 n329__vddio vss 71.1738e-18
c2022 n332__vddio vss 31.5657e-18
c2023 n333__vddio vss 29.1759e-18
c2024 n336__vddio vss 19.9241e-18
c2025 n448__i18__net5 vss 9.30995e-18
c2026 n22__reset vss 298.658e-18
c2027 n535__r_out vss 3.11627e-18
c2028 n536__r_out vss 5.90675e-18
c2029 n447__i18__net5 vss 9.30995e-18
c2030 n9__i14__net3 vss 19.7574e-18
c2031 n12__i14__net3 vss 19.4164e-18
c2032 n13__i14__net3 vss 514.824e-18
c2033 n16__i14__net3 vss 515.217e-18
c2034 n321__vddio vss 63.4059e-18
c2035 n324__vddio vss 28.7984e-18
c2036 n325__vddio vss 26.0752e-18
c2037 n328__vddio vss 17.3818e-18
c2038 n439__i18__net5 vss 9.30995e-18
c2039 n513__r_out vss 2.06465e-18
c2040 n516__r_out vss 6.75182e-18
c2041 n39__i14__net10 vss 255.42e-18
c2042 n43__i14__net10 vss 238.59e-18
c2043 n433__i18__net5 vss 9.30995e-18
c2044 n8__i14__i17__net7 vss 133.435e-18
c2045 n23__i14__net9 vss 290.044e-18
c2046 n27__i14__net9 vss 270.146e-18
c2047 n313__vddio vss 67.1012e-18
c2048 n316__vddio vss 30.1531e-18
c2049 n317__vddio vss 27.5452e-18
c2050 n320__vddio vss 18.8388e-18
c2051 n13__i14__i17__net1 vss 109.549e-18
c2052 n432__i18__net5 vss 9.41857e-18
c2053 n8__i14__i17__net1 vss 467.652e-18
c2054 n9__i14__i17__net1 vss 121.722e-18
c2055 n5__i14__i17__net8 vss 155.883e-18
c2056 n4__i14__i17__net8 vss 533.342e-18
c2057 n500__r_out vss 3.47703e-18
c2058 n503__r_out vss 6.88348e-18
c2059 n8__i14__i17__net6 vss 772.141e-18
c2060 n9__i14__i17__net6 vss 785.428e-18
c2061 n427__i18__net5 vss 9.41857e-18
c2062 n14__reset vss 433.57e-18
c2063 n15__reset vss 430.32e-18
c2064 n305__vddio vss 69.7974e-18
c2065 n308__vddio vss 31.1398e-18
c2066 n309__vddio vss 28.5257e-18
c2067 n312__vddio vss 19.5952e-18
c2068 n12__reset vss 26.2837e-18
c2069 n422__i18__net5 vss 9.20133e-18
c2070 n4__x3 vss 120.391e-18
c2071 n4__x2 vss 114.585e-18
c2072 n488__r_out vss 8.92661e-18
c2073 n417__i18__net5 vss 9.20133e-18
c2074 n297__vddio vss 68.3976e-18
c2075 n300__vddio vss 30.313e-18
c2076 n301__vddio vss 27.6064e-18
c2077 n304__vddio vss 18.6523e-18
c2078 n412__i18__net5 vss 9.30995e-18
c2079 n475__r_out vss 7.99572e-18
c2080 n404__i18__net5 vss 9.30995e-18
c2081 n289__vddio vss 66.3658e-18
c2082 n292__vddio vss 29.3337e-18
c2083 n293__vddio vss 26.7873e-18
c2084 n296__vddio vss 18.0374e-18
c2085 n401__i18__net5 vss 9.30995e-18
c2086 n470__r_out vss 9.4276e-18
c2087 n394__i18__net5 vss 9.30995e-18
c2088 n281__vddio vss 67.4376e-18
c2089 n284__vddio vss 30.1538e-18
c2090 n285__vddio vss 27.6986e-18
c2091 n288__vddio vss 18.9925e-18
c2092 n389__i18__net5 vss 9.30995e-18
c2093 n454__r_out vss 8.07667e-18
c2094 n384__i18__net5 vss 9.41857e-18
c2095 n273__vddio vss 72.2798e-18
c2096 n276__vddio vss 32.4552e-18
c2097 n277__vddio vss 30.2336e-18
c2098 n280__vddio vss 21.0047e-18
c2099 n382__i18__net5 vss 9.41857e-18
c2100 n433__r_out vss 9.55644e-18
c2101 n374__i18__net5 vss 9.20133e-18
c2102 n265__vddio vss 72.0197e-18
c2103 n268__vddio vss 31.5657e-18
c2104 n269__vddio vss 29.1759e-18
c2105 n272__vddio vss 19.9241e-18
c2106 n372__i18__net5 vss 9.20133e-18
c2107 n426__r_out vss 8.91582e-18
c2108 n364__i18__net5 vss 9.30995e-18
c2109 n257__vddio vss 65.7526e-18
c2110 n260__vddio vss 28.7984e-18
c2111 n261__vddio vss 26.0752e-18
c2112 n264__vddio vss 17.3818e-18
c2113 n359__i18__net5 vss 9.30995e-18
c2114 n413__r_out vss 8.01951e-18
c2115 n354__i18__net5 vss 9.30995e-18
c2116 n249__vddio vss 67.4302e-18
c2117 n252__vddio vss 30.3175e-18
c2118 n253__vddio vss 27.6831e-18
c2119 n256__vddio vss 18.9393e-18
c2120 n352__i18__net5 vss 9.30995e-18
c2121 n392__r_out vss 9.31657e-18
c2122 n344__i18__net5 vss 9.30995e-18
c2123 n241__vddio vss 68.7287e-18
c2124 n244__vddio vss 30.313e-18
c2125 n245__vddio vss 27.6064e-18
c2126 n248__vddio vss 18.6696e-18
c2127 n342__i18__net5 vss 9.30995e-18
c2128 n379__r_out vss 8.0309e-18
c2129 n334__i18__net5 vss 9.41857e-18
c2130 n233__vddio vss 66.3658e-18
c2131 n236__vddio vss 29.3337e-18
c2132 n237__vddio vss 26.7873e-18
c2133 n240__vddio vss 18.1527e-18
c2134 n332__i18__net5 vss 9.41857e-18
c2135 n366__r_out vss 9.56009e-18
c2136 n324__i18__net5 vss 9.20133e-18
c2137 n225__vddio vss 67.8399e-18
c2138 n228__vddio vss 30.1538e-18
c2139 n229__vddio vss 27.6986e-18
c2140 n232__vddio vss 18.9925e-18
c2141 n319__i18__net5 vss 9.20133e-18
c2142 n353__r_out vss 8.93037e-18
c2143 n317__i18__net5 vss 9.30995e-18
c2144 n217__vddio vss 72.5217e-18
c2145 n220__vddio vss 32.4552e-18
c2146 n221__vddio vss 30.2336e-18
c2147 n224__vddio vss 21.045e-18
c2148 n309__i18__net5 vss 9.30995e-18
c2149 n348__r_out vss 8.03048e-18
c2150 n307__i18__net5 vss 9.30995e-18
c2151 n209__vddio vss 71.4257e-18
c2152 n212__vddio vss 31.5657e-18
c2153 n213__vddio vss 29.1759e-18
c2154 n216__vddio vss 19.9241e-18
c2155 n302__i18__net5 vss 9.30995e-18
c2156 n327__r_out vss 9.3289e-18
c2157 n297__i18__net5 vss 9.30995e-18
c2158 n201__vddio vss 65.8596e-18
c2159 n204__vddio vss 28.7984e-18
c2160 n205__vddio vss 26.0752e-18
c2161 n208__vddio vss 17.3818e-18
c2162 n292__i18__net5 vss 9.30995e-18
c2163 n314__r_out vss 8.03493e-18
c2164 n287__i18__net5 vss 9.41857e-18
c2165 n193__vddio vss 67.1152e-18
c2166 n196__vddio vss 30.1531e-18
c2167 n197__vddio vss 27.5452e-18
c2168 n200__vddio vss 18.8388e-18
c2169 n282__i18__net5 vss 9.41857e-18
c2170 n301__r_out vss 9.55644e-18
c2171 n274__i18__net5 vss 9.20133e-18
c2172 n185__vddio vss 69.767e-18
c2173 n188__vddio vss 31.1398e-18
c2174 n189__vddio vss 28.5257e-18
c2175 n192__vddio vss 19.5952e-18
c2176 n272__i18__net5 vss 9.20133e-18
c2177 n288__r_out vss 8.91808e-18
c2178 n264__i18__net5 vss 9.30995e-18
c2179 n177__vddio vss 68.414e-18
c2180 n180__vddio vss 30.313e-18
c2181 n181__vddio vss 27.6064e-18
c2182 n184__vddio vss 18.6915e-18
c2183 n262__i18__net5 vss 9.30995e-18
c2184 n283__r_out vss 8.01951e-18
c2185 n257__i18__net5 vss 9.30995e-18
c2186 n169__vddio vss 66.3797e-18
c2187 n172__vddio vss 29.3337e-18
c2188 n173__vddio vss 26.7873e-18
c2189 n176__vddio vss 18.075e-18
c2190 n249__i18__net5 vss 9.30995e-18
c2191 n262__r_out vss 9.32383e-18
c2192 n244__i18__net5 vss 9.30995e-18
c2193 n161__vddio vss 67.5903e-18
c2194 n164__vddio vss 30.1538e-18
c2195 n165__vddio vss 27.6986e-18
c2196 n168__vddio vss 19.0042e-18
c2197 n239__i18__net5 vss 9.41857e-18
c2198 n249__r_out vss 8.02761e-18
c2199 n234__i18__net5 vss 9.41857e-18
c2200 n153__vddio vss 83.3612e-18
c2201 n156__vddio vss 43.5077e-18
c2202 n157__vddio vss 30.2336e-18
c2203 n160__vddio vss 21.0052e-18
c2204 n232__i18__net5 vss 9.20133e-18
c2205 n236__r_out vss 9.55644e-18
c2206 n227__i18__net5 vss 9.20133e-18
c2207 n145__vddio vss 68.5054e-18
c2208 n148__vddio vss 36.1171e-18
c2209 n149__vddio vss 29.1759e-18
c2210 n152__vddio vss 19.9241e-18
c2211 n222__i18__net5 vss 9.30995e-18
c2212 n223__r_out vss 8.91582e-18
c2213 n217__i18__net5 vss 9.30995e-18
c2214 n137__vddio vss 62.2026e-18
c2215 n140__vddio vss 33.3443e-18
c2216 n141__vddio vss 26.0752e-18
c2217 n144__vddio vss 17.3818e-18
c2218 n212__i18__net5 vss 9.30995e-18
c2219 n218__r_out vss 8.01951e-18
c2220 n207__i18__net5 vss 9.30995e-18
c2221 n129__vddio vss 63.0095e-18
c2222 n132__vddio vss 34.213e-18
c2223 n133__vddio vss 27.1317e-18
c2224 n136__vddio vss 18.5375e-18
c2225 n202__i18__net5 vss 9.30995e-18
c2226 n197__r_out vss 9.65225e-18
c2227 n197__i18__net5 vss 9.30995e-18
c2228 n121__vddio vss 63.2859e-18
c2229 n124__vddio vss 35.0351e-18
c2230 n125__vddio vss 27.9697e-18
c2231 n128__vddio vss 19.1888e-18
c2232 n192__i18__net5 vss 10.8719e-18
c2233 n184__r_out vss 8.0309e-18
c2234 n184__i18__net5 vss 21.2126e-18
c2235 n113__vddio vss 65.1597e-18
c2236 n116__vddio vss 34.7062e-18
c2237 n117__vddio vss 27.5382e-18
c2238 n120__vddio vss 18.8318e-18
c2239 n182__i18__net5 vss 13.9479e-18
c2240 n171__r_out vss 9.19685e-18
c2241 n177__i18__net5 vss 9.20133e-18
c2242 n105__vddio vss 63.149e-18
c2243 n108__vddio vss 33.3351e-18
c2244 n109__vddio vss 26.0543e-18
c2245 n112__vddio vss 17.4746e-18
c2246 n169__i18__net5 vss 9.47726e-18
c2247 n158__r_out vss 8.92812e-18
c2248 n167__i18__net5 vss 9.30995e-18
c2249 n97__vddio vss 67.2421e-18
c2250 n100__vddio vss 35.59e-18
c2251 n101__vddio vss 28.6575e-18
c2252 n104__vddio vss 19.3827e-18
c2253 n159__i18__net5 vss 9.30995e-18
c2254 n153__r_out vss 8.03048e-18
c2255 n157__i18__net5 vss 9.30995e-18
c2256 n89__vddio vss 68e-18
c2257 n92__vddio vss 36.1261e-18
c2258 n93__vddio vss 29.2381e-18
c2259 n96__vddio vss 20.0031e-18
c2260 n152__i18__net5 vss 9.30995e-18
c2261 n140__r_out vss 9.33114e-18
c2262 n147__i18__net5 vss 9.30995e-18
c2263 n81__vddio vss 67.4377e-18
c2264 n84__vddio vss 34.7799e-18
c2265 n85__vddio vss 26.7873e-18
c2266 n88__vddio vss 18.0744e-18
c2267 n142__i18__net5 vss 9.41857e-18
c2268 n119__r_out vss 8.03493e-18
c2269 n134__i18__net5 vss 9.41857e-18
c2270 n73__vddio vss 67.2508e-18
c2271 n76__vddio vss 30.1538e-18
c2272 n77__vddio vss 27.6986e-18
c2273 n80__vddio vss 18.9925e-18
c2274 n132__i18__net5 vss 9.20133e-18
c2275 n106__r_out vss 9.55644e-18
c2276 n127__i18__net5 vss 9.20133e-18
c2277 n65__vddio vss 61.5342e-18
c2278 n68__vddio vss 26.9659e-18
c2279 n69__vddio vss 26.2798e-18
c2280 n72__vddio vss 19.5944e-18
c2281 n118__i18__net5 vss 9.30995e-18
c2282 n93__r_out vss 8.91808e-18
c2283 n114__i18__net5 vss 9.30995e-18
c2284 n57__vddio vss 58.2027e-18
c2285 n60__vddio vss 22.8671e-18
c2286 n61__vddio vss 24.0669e-18
c2287 n64__vddio vss 19.5889e-18
c2288 n108__i18__net5 vss 9.30995e-18
c2289 n88__r_out vss 8.01951e-18
c2290 n107__i18__net5 vss 9.30995e-18
c2291 n49__vddio vss 56.338e-18
c2292 n52__vddio vss 22.111e-18
c2293 n53__vddio vss 23.1997e-18
c2294 n56__vddio vss 18.8304e-18
c2295 n99__i18__net5 vss 9.30995e-18
c2296 n67__r_out vss 9.31657e-18
c2297 n94__i18__net5 vss 9.41857e-18
c2298 n41__vddio vss 55.718e-18
c2299 n44__vddio vss 20.7426e-18
c2300 n45__vddio vss 21.7189e-18
c2301 n48__vddio vss 17.2419e-18
c2302 n89__i18__net5 vss 9.41857e-18
c2303 n54__r_out vss 8.02864e-18
c2304 n84__i18__net5 vss 9.20133e-18
c2305 n33__vddio vss 59.4782e-18
c2306 n36__vddio vss 22.4588e-18
c2307 n37__vddio vss 24.0496e-18
c2308 n40__vddio vss 19.4185e-18
c2309 n82__i18__net5 vss 9.20133e-18
c2310 n41__r_out vss 9.56009e-18
c2311 n77__i18__net5 vss 9.30995e-18
c2312 n25__vddio vss 60.8055e-18
c2313 n28__vddio vss 22.9949e-18
c2314 n29__vddio vss 24.6302e-18
c2315 n32__vddio vss 20.0411e-18
c2316 n72__i18__net5 vss 9.30995e-18
c2317 n28__r_out vss 8.93037e-18
c2318 n67__i18__net5 vss 9.30995e-18
c2319 n17__vddio vss 55.4945e-18
c2320 n20__vddio vss 21.291e-18
c2321 n21__vddio vss 22.4488e-18
c2322 n24__vddio vss 18.0735e-18
c2323 n59__i18__net5 vss 9.30995e-18
c2324 n23__r_out vss 8.04017e-18
c2325 n57__i18__net5 vss 9.30995e-18
c2326 n9__vddio vss 56.5224e-18
c2327 n12__vddio vss 22.1111e-18
c2328 n13__vddio vss 23.36e-18
c2329 n16__vddio vss 18.991e-18
c2330 n49__i18__net5 vss 9.76304e-18
c2331 n2__r_out vss 12.2504e-18
c2332 n47__i18__net5 vss 19.6675e-18
c2333 n1__vddio vss 36.2983e-18
c2334 n4__vddio vss 11.7889e-18
c2335 n5__vddio vss 12.9758e-18
c2336 n8__vddio vss 10.6706e-18
c2337 n8__serial_out_b_high_buff vss 290.136e-18
c2338 n4__serial_out_b_high_buff vss 372.016e-18
c2339 n12__r0_buff vss 33.8282e-18
c2340 n10__r2_buff vss 33.0543e-18
c2341 n12__r1_buff vss 35.3565e-18
c2342 n684__vddio vss 52.7625e-18
c2343 n670__vddio vss 75.4774e-18
c2344 n13__serial_out_b_high vss 36.3269e-18
c2345 n31__vdd vss 214.555e-18
c2346 n131__vdd vss 152.016e-18
c2347 n24__serial_out vss 113.239e-18
c2348 n680__vddio vss 23.458e-18
c2349 n9__r2 vss 26.7654e-18
c2350 n14__r0 vss 16.4338e-18
c2351 n13__r1 vss 19.1485e-18
c2352 n12__serial_out_b_high vss 76.6705e-18
c2353 n661__vddio vss 26.9346e-18
c2354 n8__i12__bio vss 247.426e-18
c2355 n2__i2__q vss 126.569e-18
c2356 n2__i1__q vss 146.425e-18
c2357 n2__i0__q vss 168.097e-18
c2358 n11__serial_out_b_high vss 140.863e-18
c2359 n22__serial_out vss 51.2472e-18
c2360 n13__net4 vss 54.729e-18
c2361 n12__net3 vss 48.4848e-18
c2362 n4__i12__bio vss 165.262e-18
c2363 n13__i2__net77 vss 89.8253e-18
c2364 n13__i1__net77 vss 91.2794e-18
c2365 n13__i0__net77 vss 89.3112e-18
c2366 n7__i12__bio vss 186.452e-18
c2367 n7__serial_out_b_high vss 117.629e-18
c2368 n9__i2__net77 vss 78.6975e-18
c2369 n9__i1__net77 vss 81.7681e-18
c2370 n9__i0__net77 vss 76.5357e-18
c2371 n12__i2__net77 vss 92.547e-18
c2372 n12__i1__net77 vss 121.395e-18
c2373 n12__i0__net77 vss 121.499e-18
c2374 n14__i2__net76 vss 143.071e-18
c2375 n14__i1__net76 vss 151.661e-18
c2376 n14__i0__net76 vss 143.969e-18
c2377 n25__reset_b vss 304.718e-18
c2378 n26__reset_b vss 298.609e-18
c2379 n27__reset_b vss 314.384e-18
c2380 n639__vddio vss 12.7528e-18
c2381 n12__r1 vss 116.658e-18
c2382 n49__i18__net3 vss 59.5174e-18
c2383 n7__i2__net77 vss 141.318e-18
c2384 n7__i1__net77 vss 158.076e-18
c2385 n7__i0__net77 vss 159.084e-18
c2386 n7__i13__i20__i4__net2 vss 61.6294e-18
c2387 n27__i13__net18 vss 70.3743e-18
c2388 n198__i18__net4 vss 61.1236e-18
c2389 n201__i18__net4 vss 72.8469e-18
c2390 n20__i13__net7 vss 131.913e-18
c2391 n11__i2__net76 vss 116.295e-18
c2392 n11__i1__net76 vss 122.829e-18
c2393 n11__i0__net76 vss 112.843e-18
c2394 n46__i18__net3 vss 61.12e-21
c2395 n8__r1 vss 432.238e-18
c2396 n6__i13__i20__i4__net2 vss 137.166e-18
c2397 n44__ck_b vss 178.996e-18
c2398 n47__ck_buff vss 202.773e-18
c2399 n48__ck_buff vss 251.379e-18
c2400 n45__ck_b vss 177.092e-18
c2401 n46__ck_b vss 177.576e-18
c2402 n49__ck_buff vss 199.393e-18
c2403 n23__i13__net18 vss 133.049e-18
c2404 n642__vddio vss 48.298e-18
c2405 n17__i13__net7 vss 138.159e-18
c2406 n45__i18__net3 vss 61.12e-21
c2407 n24__i13__net18 vss 199.032e-18
c2408 n187__i18__net4 vss 58.5197e-18
c2409 n190__i18__net4 vss 71.1839e-18
c2410 n4__i13__i20__i4__net2 vss 134.887e-18
c2411 n43__i18__net3 vss 61.12e-21
c2412 n22__i13__net18 vss 193.145e-18
c2413 n5__i2__net75 vss 197.208e-18
c2414 n5__i1__net75 vss 217.139e-18
c2415 n5__i0__net75 vss 216.732e-18
c2416 n41__i18__net3 vss 61.12e-21
c2417 n6__i13__net23 vss 34.3819e-18
c2418 n2__r2 vss 85.2155e-18
c2419 n16__i2__net74 vss 118.729e-18
c2420 n16__i1__net74 vss 136.339e-18
c2421 n16__i0__net74 vss 126.271e-18
c2422 n178__i18__net4 vss 64.5389e-18
c2423 n179__i18__net4 vss 71.2505e-18
c2424 n30__reset_buff vss 444.91e-18
c2425 n31__reset_buff vss 495.634e-18
c2426 n32__reset_buff vss 440.692e-18
c2427 n39__i18__net3 vss 61.12e-21
c2428 n15__i2__net74 vss 268.077e-18
c2429 n15__i1__net74 vss 303.009e-18
c2430 n15__i0__net74 vss 266.951e-18
c2431 n41__ck_b vss 341.349e-18
c2432 n42__ck_b vss 348.027e-18
c2433 n43__ck_b vss 349.529e-18
c2434 n7__i13__i20__net1 vss 37.8429e-18
c2435 n6__i13__net3 vss 42.9178e-18
c2436 n36__i18__net3 vss 61.12e-21
c2437 n5__i13__net23 vss 148.688e-18
c2438 n20__i13__net18 vss 189.882e-18
c2439 n41__ck_buff vss 244.517e-18
c2440 n42__ck_buff vss 283.18e-18
c2441 n43__ck_buff vss 300.361e-18
c2442 n44__ck_buff vss 246.438e-18
c2443 n45__ck_buff vss 245.855e-18
c2444 n46__ck_buff vss 286.978e-18
c2445 n165__i18__net4 vss 65.526e-18
c2446 n168__i18__net4 vss 71.2434e-18
c2447 n9__i13__net17 vss 126.993e-18
c2448 n5__i13__i20__net1 vss 105.147e-18
c2449 n5__i13__net3 vss 115.377e-18
c2450 n14__i13__net7 vss 207.455e-18
c2451 n38__ck_b vss 277.761e-18
c2452 n39__ck_b vss 283.544e-18
c2453 n40__ck_b vss 281.453e-18
c2454 n35__i18__net3 vss 61.12e-21
c2455 n4__i2__net75 vss 228.214e-18
c2456 n4__i1__net75 vss 248.51e-18
c2457 n4__i0__net75 vss 249.68e-18
c2458 n33__i18__net3 vss 546.064e-21
c2459 n11__i2__net74 vss 220.857e-18
c2460 n11__i1__net74 vss 251.154e-18
c2461 n11__i0__net74 vss 229.04e-18
c2462 n154__i18__net4 vss 59.5722e-18
c2463 n157__i18__net4 vss 80.7015e-18
c2464 n38__ck_buff vss 213.938e-18
c2465 n35__ck_b vss 318.288e-18
c2466 n36__ck_b vss 360.705e-18
c2467 n39__ck_buff vss 224.155e-18
c2468 n40__ck_buff vss 223.692e-18
c2469 n37__ck_b vss 328.028e-18
c2470 n31__i18__net3 vss 6.51734e-18
c2471 n18__i13__net18 vss 80.3768e-18
c2472 n7__r0 vss 68.9365e-18
c2473 n7__i13__i19__i4__net2 vss 91.6965e-18
c2474 n23__i13__net1 vss 70.3204e-18
c2475 n27__i13__net2 vss 69.824e-18
c2476 n10__i13__i18__i4__net2 vss 116.089e-18
c2477 n20__i13__net11 vss 133.003e-18
c2478 n24__i13__net12 vss 128.991e-18
c2479 n14__i13__net18 vss 194.398e-18
c2480 n4__r0 vss 194.249e-18
c2481 n6__i13__i19__i4__net2 vss 136.724e-18
c2482 n6__i13__i18__i4__net2 vss 134.546e-18
c2483 n21__i13__net1 vss 134.217e-18
c2484 n25__i13__net2 vss 134.195e-18
c2485 n17__i13__net11 vss 136.969e-18
c2486 n21__i13__net12 vss 136.452e-18
c2487 n19__i13__net1 vss 196.509e-18
c2488 n23__i13__net2 vss 195.854e-18
c2489 n4__i13__i19__i4__net2 vss 133.273e-18
c2490 n4__i13__i18__i4__net2 vss 145.943e-18
c2491 n537__vddio vss 83.7502e-18
c2492 n539__vddio vss 81.6646e-18
c2493 n541__vddio vss 61.2722e-18
c2494 n543__vddio vss 47.5924e-18
c2495 n18__i13__net1 vss 191.777e-18
c2496 n22__i13__net2 vss 192.759e-18
c2497 n149__i18__net4 vss 29.5817e-18
c2498 n687__i18__net5 vss 69.8456e-18
c2499 n691__i18__net5 vss 70.8341e-18
c2500 n5__i13__net17 vss 256.838e-18
c2501 n9__i13__net7 vss 187.035e-18
c2502 n23__vdd vss 40.2404e-18
c2503 n147__i18__net4 vss 61.12e-21
c2504 n4__r0_buff vss 83.5333e-18
c2505 n4__r1_buff vss 84.5103e-18
c2506 n4__r2_buff vss 84.8759e-18
c2507 n529__vddio vss 142.261e-18
c2508 n532__vddio vss 128.668e-18
c2509 n533__vddio vss 76.3798e-18
c2510 n37__shift vss 174.155e-18
c2511 n38__shift vss 170.21e-18
c2512 n39__shift vss 174.409e-18
c2513 n145__i18__net4 vss 61.12e-21
c2514 n11__i2__net79 vss 147.282e-18
c2515 n11__i1__net79 vss 146.082e-18
c2516 n11__i0__net79 vss 148.984e-18
c2517 n7__i13__i19__net1 vss 35.5908e-18
c2518 n7__i13__i18__net1 vss 35.1612e-18
c2519 n672__i18__net5 vss 58.5197e-18
c2520 n673__i18__net5 vss 69.7672e-18
c2521 n34__shift vss 184.1e-18
c2522 n35__shift vss 189.499e-18
c2523 n36__shift vss 186.934e-18
c2524 n17__i13__net1 vss 190.617e-18
c2525 n21__i13__net2 vss 164.076e-18
c2526 n10__i2__net79 vss 137.882e-18
c2527 n10__i1__net79 vss 163.365e-18
c2528 n10__i0__net79 vss 163.858e-18
c2529 n2__net4 vss 69.2492e-18
c2530 n143__i18__net4 vss 61.12e-21
c2531 n5__i13__i19__net1 vss 104.466e-18
c2532 n6__i13__i18__net1 vss 104.365e-18
c2533 n15__i13__net11 vss 209.418e-18
c2534 n19__i13__net12 vss 226.464e-18
c2535 n5__i2__net79 vss 78.0121e-18
c2536 n5__i1__net79 vss 76.8046e-18
c2537 n5__i0__net79 vss 82.2676e-18
c2538 n8__i2__net79 vss 117.825e-18
c2539 n8__i1__net79 vss 126.457e-18
c2540 n8__i0__net79 vss 124.841e-18
c2541 n523__vddio vss 144.669e-18
c2542 n526__vddio vss 131.641e-18
c2543 n527__vddio vss 79.3173e-18
c2544 n31__shift vss 96.8277e-18
c2545 n32__shift vss 95.8035e-18
c2546 n33__shift vss 190.243e-18
c2547 n141__i18__net4 vss 61.12e-21
c2548 n661__i18__net5 vss 58.7858e-18
c2549 n665__i18__net5 vss 76.6627e-18
c2550 n139__i18__net4 vss 61.12e-21
c2551 n5__i9__i1__net1 vss 89.1815e-18
c2552 n517__vddio vss 143.265e-18
c2553 n520__vddio vss 131.641e-18
c2554 n521__vddio vss 78.5847e-18
c2555 n30__shift vss 85.513e-18
c2556 n548__vddio vss 52.5434e-18
c2557 n137__i18__net4 vss 61.12e-21
c2558 n16__i13__net12 vss 80.6063e-18
c2559 n17__i13__net2 vss 90.4724e-18
c2560 n16__ck4 vss 106.098e-18
c2561 n4__i9__i1__net1 vss 102.647e-18
c2562 n648__i18__net5 vss 65.5426e-18
c2563 n652__i18__net5 vss 69.827e-18
c2564 n7__i13__i17__i4__net2 vss 51.6756e-18
c2565 n29__i13__a2 vss 73.7554e-18
c2566 n29__i13__a0 vss 73.6911e-18
c2567 n10__i13__i16__i4__net2 vss 46.3471e-18
c2568 n24__i13__a3 vss 131.951e-18
c2569 n24__i13__a1 vss 131.15e-18
c2570 n14__reset_buff vss 84.3874e-18
c2571 n135__i18__net4 vss 61.12e-21
c2572 n26__shift vss 72.1704e-18
c2573 n28__shift vss 109.91e-18
c2574 n12__i13__net12 vss 194.429e-18
c2575 n14__i13__net2 vss 194.564e-18
c2576 n15__net14 vss 126.179e-18
c2577 n10__i9__net1 vss 82.9186e-18
c2578 n2__i9__i1__net1 vss 73.0725e-18
c2579 n511__vddio vss 143.762e-18
c2580 n514__vddio vss 131.641e-18
c2581 n515__vddio vss 78.5847e-18
c2582 n6__i13__i17__i4__net2 vss 135.067e-18
c2583 n6__i13__i16__i4__net2 vss 134.232e-18
c2584 n27__i13__a2 vss 134.231e-18
c2585 n27__i13__a0 vss 134.254e-18
c2586 n133__i18__net4 vss 61.12e-21
c2587 n21__i13__a3 vss 135.591e-18
c2588 n21__i13__a1 vss 135.585e-18
c2589 n11__reset_buff vss 102.935e-18
c2590 n25__i13__a2 vss 195.334e-18
c2591 n25__i13__a0 vss 194.994e-18
c2592 n636__i18__net5 vss 64.313e-18
c2593 n637__i18__net5 vss 69.7672e-18
c2594 n14__net14 vss 101.057e-18
c2595 n4__i13__i17__i4__net2 vss 131.829e-18
c2596 n4__i13__i16__i4__net2 vss 145.82e-18
c2597 n8__i9__net1 vss 110.092e-18
c2598 n131__i18__net4 vss 61.12e-21
c2599 n25__ck_buff vss 48.4905e-18
c2600 n24__i13__a2 vss 188.964e-18
c2601 n24__i13__a0 vss 187.418e-18
c2602 n15__net13 vss 114.606e-18
c2603 n506__vddio vss 135.809e-18
c2604 n507__vddio vss 137.149e-18
c2605 n510__vddio vss 73.0091e-18
c2606 n129__i18__net4 vss 61.12e-21
c2607 n7__i9__net2 vss 104.024e-18
c2608 n63__reset vss 73.4383e-18
c2609 n9__i13__net11 vss 205.757e-18
c2610 n11__i13__net1 vss 151.583e-18
c2611 n14__ck_buff vss 108.385e-18
c2612 n622__i18__net5 vss 199.73e-18
c2613 n626__i18__net5 vss 76.8208e-18
c2614 n13__i9__i4__net4 vss 88.3779e-18
c2615 n11__net13 vss 89.2331e-18
c2616 n127__i18__net4 vss 61.12e-21
c2617 n60__reset vss 28.9221e-18
c2618 n500__vddio vss 141.694e-18
c2619 n501__vddio vss 129.703e-18
c2620 n504__vddio vss 71.3477e-18
c2621 n7__i13__i17__net1 vss 34.8081e-18
c2622 n7__i13__i16__net1 vss 34.3946e-18
c2623 n9__i9__i4__net4 vss 72.5804e-18
c2624 n125__i18__net4 vss 61.12e-21
c2625 n12__i9__i4__net4 vss 116.682e-18
c2626 n23__i13__a2 vss 181.168e-18
c2627 n23__i13__a0 vss 162.345e-18
c2628 n609__i18__net5 vss 64.368e-18
c2629 n613__i18__net5 vss 69.8309e-18
c2630 n5__i13__i17__net1 vss 107.85e-18
c2631 n6__i13__i16__net1 vss 108.269e-18
c2632 n19__i13__a3 vss 201.187e-18
c2633 n19__i13__a1 vss 201.055e-18
c2634 n123__i18__net4 vss 61.12e-21
c2635 n34__ck vss 74.3163e-18
c2636 n14__i9__i4__net5 vss 144.877e-18
c2637 n493__vddio vss 142.888e-18
c2638 n496__vddio vss 129.703e-18
c2639 n497__vddio vss 77.7863e-18
c2640 n14__reset_b vss 205.143e-18
c2641 n553__vddio vss 52.3011e-18
c2642 n119__i18__net4 vss 61.12e-21
c2643 n593__i18__net5 vss 125.789e-18
c2644 n596__i18__net5 vss 76.5972e-18
c2645 n116__i18__net4 vss 61.12e-21
c2646 n7__i9__i4__net4 vss 150.401e-18
c2647 n16__i13__a3 vss 89.0926e-18
c2648 n15__i13__a1 vss 88.7463e-18
c2649 n487__vddio vss 46.2528e-18
c2650 n490__vddio vss 37.4346e-18
c2651 n491__vddio vss 43.9487e-18
c2652 n11__i9__i4__net5 vss 120.737e-18
c2653 n108__i18__net4 vss 61.12e-21
c2654 n12__net12 vss 84.2435e-18
c2655 n7__i13__i15__net2 vss 28.3665e-18
c2656 n22__x_out_3 vss 76.0211e-18
c2657 n23__x_out_1 vss 75.4144e-18
c2658 n10__i13__i13__net2 vss 29.2955e-18
c2659 n583__i18__net5 vss 209.096e-18
c2660 n587__i18__net5 vss 69.7478e-18
c2661 n18__y_out_3 vss 133.396e-18
c2662 n19__y_out_1 vss 133.828e-18
c2663 n18__ck_b vss 183.822e-18
c2664 n12__ck_buff vss 204.987e-18
c2665 n11__reset_b vss 109.771e-18
c2666 n12__i13__a3 vss 201.089e-18
c2667 n12__i13__a1 vss 201.425e-18
c2668 n106__i18__net4 vss 61.12e-21
c2669 n6__i13__i15__net2 vss 135.264e-18
c2670 n6__i13__i13__net2 vss 136.71e-18
c2671 n20__x_out_3 vss 141.436e-18
c2672 n19__x_out_1 vss 139.282e-18
c2673 n11__net12 vss 114.959e-18
c2674 n14__y_out_3 vss 137.741e-18
c2675 n13__y_out_1 vss 136.023e-18
c2676 n481__vddio vss 45.601e-18
c2677 n484__vddio vss 37.4346e-18
c2678 n485__vddio vss 43.2971e-18
c2679 n8__reset_b vss 115.284e-18
c2680 n98__i18__net4 vss 61.12e-21
c2681 n18__x_out_3 vss 197.568e-18
c2682 n17__x_out_1 vss 194.544e-18
c2683 n30__ck vss 91.1388e-18
c2684 n4__i13__i15__net2 vss 114.806e-18
c2685 n4__i13__i13__net2 vss 132.089e-18
c2686 n5__i9__i4__net2 vss 204.704e-18
c2687 n570__i18__net5 vss 64.0684e-18
c2688 n574__i18__net5 vss 69.8231e-18
c2689 n17__x_out_3 vss 76.3754e-18
c2690 n16__x_out_1 vss 73.5727e-18
c2691 n94__i18__net4 vss 61.12e-21
c2692 n16__i9__i4__net1 vss 114.259e-18
c2693 n475__vddio vss 142.631e-18
c2694 n478__vddio vss 131.217e-18
c2695 n479__vddio vss 77.9252e-18
c2696 n91__i18__net4 vss 61.12e-21
c2697 n14__i9__i4__net1 vss 255.793e-18
c2698 n17__ck_b vss 331.454e-18
c2699 n554__i18__net5 vss 59.3179e-18
c2700 n557__i18__net5 vss 76.8844e-18
c2701 n86__i18__net4 vss 61.12e-21
c2702 n10__ck_buff vss 114.155e-18
c2703 n11__ck_buff vss 293.707e-18
c2704 n469__vddio vss 141.049e-18
c2705 n472__vddio vss 129.703e-18
c2706 n473__vddio vss 76.6714e-18
c2707 n16__ck_b vss 274.271e-18
c2708 n18__i13__a2 vss 85.743e-18
c2709 n17__i13__a0 vss 80.6502e-18
c2710 n558__vddio vss 52.5634e-18
c2711 n78__i18__net4 vss 61.12e-21
c2712 n7__i13__i14__net2 vss 32.6091e-18
c2713 n23__x_out_2 vss 73.8286e-18
c2714 n19__y_out_0 vss 73.3651e-18
c2715 n10__i13__i12__net2 vss 29.9642e-18
c2716 n544__i18__net5 vss 58.2537e-18
c2717 n548__i18__net5 vss 69.7672e-18
c2718 n4__i9__i4__net2 vss 243.899e-18
c2719 n19__y_out_2 vss 125.755e-18
c2720 n19__x_out_0 vss 125.875e-18
c2721 n76__i18__net4 vss 61.12e-21
c2722 n12__i13__a2 vss 195.316e-18
c2723 n12__i13__a0 vss 194.767e-18
c2724 n12__net11 vss 87.4326e-18
c2725 n11__i9__i4__net1 vss 245.949e-18
c2726 n463__vddio vss 142.953e-18
c2727 n466__vddio vss 129.703e-18
c2728 n467__vddio vss 77.732e-18
c2729 n6__i13__i14__net2 vss 136.801e-18
c2730 n6__i13__i12__net2 vss 135.222e-18
c2731 n21__x_out_2 vss 141.708e-18
c2732 n17__y_out_0 vss 139.136e-18
c2733 n13__y_out_2 vss 136.022e-18
c2734 n15__x_out_0 vss 136.561e-18
c2735 n10__ck_b vss 88.9971e-18
c2736 n7__ck_buff vss 175.714e-18
c2737 n8__ck_b vss 313.932e-18
c2738 n71__i18__net4 vss 61.12e-21
c2739 n17__x_out_2 vss 197.49e-18
c2740 n15__y_out_0 vss 196.968e-18
c2741 n7__ck4 vss 84.1902e-18
c2742 n4__i13__i14__net2 vss 110.582e-18
c2743 n4__i13__i12__net2 vss 132.463e-18
c2744 n531__i18__net5 vss 64.2683e-18
c2745 n535__i18__net5 vss 69.8341e-18
c2746 n11__net11 vss 116.231e-18
c2747 n66__i18__net4 vss 61.12e-21
c2748 n16__x_out_2 vss 83.1871e-18
c2749 n14__y_out_0 vss 71.5909e-18
c2750 n6__ck_b vss 69.2199e-18
c2751 n458__vddio vss 133.164e-18
c2752 n459__vddio vss 135.657e-18
c2753 n462__vddio vss 70.9494e-18
c2754 n58__i18__net4 vss 61.12e-21
c2755 n8__y_out_3 vss 58.9838e-18
c2756 n8__y_out_2 vss 56.9827e-18
c2757 n8__y_out_1 vss 68.1044e-18
c2758 n10__y_out_0 vss 50.5265e-18
c2759 n518__i18__net5 vss 65.2494e-18
c2760 n522__i18__net5 vss 69.827e-18
c2761 n93__i14__net9 vss 102.485e-18
c2762 n104__i14__net10 vss 30.5352e-18
c2763 n56__i18__net4 vss 409.461e-21
c2764 n37__i14__net7 vss 116.362e-18
c2765 n36__i14__net11 vss 107.329e-18
c2766 n452__vddio vss 134.582e-18
c2767 n453__vddio vss 135.626e-18
c2768 n456__vddio vss 71.4551e-18
c2769 n8__i14__x_out_b_1 vss 292.12e-18
c2770 n9__i14__y_out_b_2 vss 291.607e-18
c2771 n8__i14__y_out_b_1 vss 294.894e-18
c2772 n9__i14__x_out_b_0 vss 298.47e-18
c2773 n51__i18__net4 vss 473.324e-21
c2774 n90__i14__net9 vss 124.31e-18
c2775 n101__i14__net10 vss 46.9506e-18
c2776 n13__i14__i11__net4 vss 91.1629e-18
c2777 n13__i14__i14__net4 vss 97.9053e-18
c2778 n13__i14__i15__net4 vss 85.5515e-18
c2779 n13__i14__i12__net4 vss 87.1487e-18
c2780 n502__i18__net5 vss 59.3013e-18
c2781 n505__i18__net5 vss 79.3752e-18
c2782 n34__i14__net7 vss 72.5246e-18
c2783 n34__i14__net11 vss 106.95e-18
c2784 n43__i18__net4 vss 6.2383e-18
c2785 n87__i14__net9 vss 116.468e-18
c2786 n98__i14__net10 vss 31.6376e-18
c2787 n10__i14__i11__net4 vss 74.7921e-18
c2788 n10__i14__i14__net4 vss 81.4805e-18
c2789 n10__i14__i15__net4 vss 70.0519e-18
c2790 n10__i14__i12__net4 vss 69.9306e-18
c2791 n429__vddio vss 83.8677e-18
c2792 n432__vddio vss 71.211e-18
c2793 n433__vddio vss 60.6632e-18
c2794 n8__i14__i11__net4 vss 109.586e-18
c2795 n8__i14__i14__net4 vss 110.158e-18
c2796 n8__i14__i15__net4 vss 109.76e-18
c2797 n8__i14__i12__net4 vss 109.946e-18
c2798 n4__ck4 vss 140.573e-18
c2799 n14__i14__i11__net5 vss 143.398e-18
c2800 n14__i14__i14__net5 vss 143.105e-18
c2801 n14__i14__i15__net5 vss 142.838e-18
c2802 n14__i14__i12__net5 vss 142.801e-18
c2803 n68__i14__net3 vss 22.5069e-18
c2804 n72__i14__net4 vss 113.092e-18
c2805 n73__i14__net4 vss 119.021e-18
c2806 n74__i14__net4 vss 107.529e-18
c2807 n75__i14__net4 vss 119.1e-18
c2808 n31__i14__net11 vss 126.033e-18
c2809 n71__i14__net4 vss 117.336e-18
c2810 n61__i14__net3 vss 35.4366e-18
c2811 n7__i14__i11__net4 vss 149.426e-18
c2812 n7__i14__i14__net4 vss 149.358e-18
c2813 n7__i14__i15__net4 vss 149.397e-18
c2814 n7__i14__i12__net4 vss 157.169e-18
c2815 n33__i14__net7 vss 79.7376e-18
c2816 n70__i14__net4 vss 119.732e-18
c2817 n29__i14__net7 vss 158.042e-18
c2818 n11__i14__i11__net5 vss 116.125e-18
c2819 n11__i14__i14__net5 vss 114.224e-18
c2820 n11__i14__i15__net5 vss 115.466e-18
c2821 n11__i14__i12__net5 vss 114.632e-18
c2822 n58__i14__net3 vss 51.5627e-18
c2823 n402__vddio vss 70.8917e-18
c2824 n403__vddio vss 66.6321e-18
c2825 n406__vddio vss 59.8964e-18
c2826 n407__vddio vss 44.4676e-18
c2827 n499__i18__net5 vss 30.796e-18
c2828 n93__i14__net10 vss 199.865e-18
c2829 n77__i14__net9 vss 177.074e-18
c2830 n78__i14__net9 vss 175.988e-18
c2831 n94__i14__net10 vss 200.236e-18
c2832 n95__i14__net10 vss 202.901e-18
c2833 n79__i14__net9 vss 177.051e-18
c2834 n80__i14__net9 vss 176.011e-18
c2835 n96__i14__net10 vss 200.393e-18
c2836 n646__r_out vss 202.241e-18
c2837 n650__r_out vss 79.6053e-18
c2838 n56__i14__net4 vss 120.115e-18
c2839 n15__i14__i17__net11 vss 139.726e-18
c2840 n497__i18__net5 vss 61.12e-21
c2841 n19__i14__i17__net10 vss 153.325e-18
c2842 n25__i14__i17__net8 vss 241.303e-18
c2843 n49__reset vss 128.836e-18
c2844 n394__vddio vss 131.382e-18
c2845 n395__vddio vss 123.983e-18
c2846 n398__vddio vss 110.605e-18
c2847 n399__vddio vss 83.9964e-18
c2848 n5__i14__i11__net2 vss 203.103e-18
c2849 n5__i14__i14__net2 vss 203.027e-18
c2850 n5__i14__i15__net2 vss 203.039e-18
c2851 n5__i14__i12__net2 vss 203.014e-18
c2852 n53__i14__net4 vss 132.217e-18
c2853 n495__i18__net5 vss 61.12e-21
c2854 n14__i14__i17__net11 vss 238.135e-18
c2855 n48__reset vss 143.104e-18
c2856 n17__i14__i17__net10 vss 143.446e-18
c2857 n633__r_out vss 64.887e-18
c2858 n637__r_out vss 78.0242e-18
c2859 n16__i14__i11__net1 vss 113.425e-18
c2860 n16__i14__i14__net1 vss 113.197e-18
c2861 n16__i14__i15__net1 vss 112.948e-18
c2862 n16__i14__i12__net1 vss 113.086e-18
c2863 n50__i14__net4 vss 112.233e-18
c2864 n38__i14__net3 vss 501.703e-18
c2865 n493__i18__net5 vss 61.12e-21
c2866 n19__i14__i17__net9 vss 260.989e-18
c2867 n14__i14__i11__net1 vss 255.112e-18
c2868 n14__i14__i14__net1 vss 254.786e-18
c2869 n14__i14__i15__net1 vss 255.05e-18
c2870 n14__i14__i12__net1 vss 254.826e-18
c2871 n385__vddio vss 139.345e-18
c2872 n388__vddio vss 117.897e-18
c2873 n389__vddio vss 116.407e-18
c2874 n392__vddio vss 89.79e-18
c2875 n12__i14__i17__net10 vss 173.545e-18
c2876 n73__i14__net9 vss 325.55e-18
c2877 n74__i14__net9 vss 325.647e-18
c2878 n75__i14__net9 vss 325.592e-18
c2879 n76__i14__net9 vss 325.21e-18
c2880 n491__i18__net5 vss 61.12e-21
c2881 n14__i14__i17__net9 vss 108.773e-18
c2882 n77__i14__net10 vss 283.525e-18
c2883 n78__i14__net10 vss 254.896e-18
c2884 n79__i14__net10 vss 254.676e-18
c2885 n80__i14__net10 vss 285.419e-18
c2886 n81__i14__net10 vss 285.222e-18
c2887 n82__i14__net10 vss 234.179e-18
c2888 n83__i14__net10 vss 234.123e-18
c2889 n84__i14__net10 vss 284.46e-18
c2890 n28__i14__net7 vss 270.811e-18
c2891 n620__r_out vss 205.161e-18
c2892 n624__r_out vss 77.2907e-18
c2893 n24__i14__i17__net8 vss 300.844e-18
c2894 n11__i14__i17__net9 vss 110.829e-18
c2895 n63__i14__net9 vss 266.207e-18
c2896 n67__i14__net9 vss 267.001e-18
c2897 n489__i18__net5 vss 61.12e-21
c2898 n13__i14__i17__net11 vss 101.559e-18
c2899 n378__vddio vss 129.727e-18
c2900 n379__vddio vss 123.522e-18
c2901 n382__vddio vss 109.373e-18
c2902 n383__vddio vss 82.4675e-18
c2903 n28__i14__net11 vss 205.083e-18
c2904 n9__i14__i17__net9 vss 140.435e-18
c2905 n4__i14__i11__net2 vss 236.097e-18
c2906 n4__i14__i14__net2 vss 236.286e-18
c2907 n4__i14__i15__net2 vss 236.286e-18
c2908 n4__i14__i12__net2 vss 235.993e-18
c2909 n487__i18__net5 vss 61.12e-21
c2910 n23__i14__i17__net8 vss 120.3e-18
c2911 n9__i14__i17__net10 vss 73.7011e-18
c2912 n11__i14__i11__net1 vss 244.44e-18
c2913 n11__i14__i14__net1 vss 243.963e-18
c2914 n11__i14__i15__net1 vss 244.148e-18
c2915 n11__i14__i12__net1 vss 244.848e-18
c2916 n607__r_out vss 205.48e-18
c2917 n611__r_out vss 85.4076e-18
c2918 n485__i18__net5 vss 61.12e-21
c2919 n66__i14__net10 vss 147.484e-18
c2920 n70__i14__net10 vss 146.612e-18
c2921 n72__i14__net10 vss 147.429e-18
c2922 n76__i14__net10 vss 146.719e-18
c2923 n18__i14__i17__net7 vss 48.5532e-18
c2924 n11__i14__i17__net11 vss 46.2061e-18
c2925 n57__i14__net9 vss 257.044e-18
c2926 n58__i14__net9 vss 254.891e-18
c2927 n59__i14__net9 vss 256.61e-18
c2928 n60__i14__net9 vss 255.363e-18
c2929 n370__vddio vss 129.729e-18
c2930 n371__vddio vss 122.806e-18
c2931 n374__vddio vss 109.373e-18
c2932 n375__vddio vss 82.4675e-18
c2933 n2__y3 vss 194.966e-18
c2934 n2__y2 vss 193.31e-18
c2935 n2__y1 vss 90.272e-18
c2936 n2__y0 vss 90.1957e-18
c2937 n483__i18__net5 vss 61.12e-21
c2938 n27__i14__i17__net1 vss 52.9429e-18
c2939 n21__i14__i17__net8 vss 33.2179e-18
c2940 n2__x_out_3 vss 83.9753e-18
c2941 n2__x_out_2 vss 81.1074e-18
c2942 n2__x_out_1 vss 46.452e-18
c2943 n2__x_out_0 vss 46.4044e-18
c2944 n594__r_out vss 64.5779e-18
c2945 n598__r_out vss 78.3286e-18
c2946 n13__i14__i17__i2__net4 vss 94.8966e-18
c2947 n13__i14__i17__i3__net4 vss 96.3154e-18
c2948 n481__i18__net5 vss 61.12e-21
c2949 n362__vddio vss 129.728e-18
c2950 n363__vddio vss 122.806e-18
c2951 n366__vddio vss 109.373e-18
c2952 n367__vddio vss 82.4675e-18
c2953 n8__i14__y_out_b_3 vss 1.79626e-15
c2954 n9__i14__y_out_b_0 vss 1.79514e-15
c2955 n8__i14__x_out_b_2 vss 1.79086e-15
c2956 n9__i14__x_out_b_3 vss 1.79201e-15
c2957 n479__i18__net5 vss 61.12e-21
c2958 n9__i14__i17__i2__net4 vss 84.2628e-18
c2959 n9__i14__i17__i3__net4 vss 79.0011e-18
c2960 n12__i14__i17__i2__net4 vss 110.382e-18
c2961 n12__i14__i17__i3__net4 vss 116.861e-18
c2962 n13__i14__i13__net4 vss 88.9485e-18
c2963 n13__i14__i16__net4 vss 89.6221e-18
c2964 n13__i14__i10__net4 vss 90.382e-18
c2965 n13__i14__i9__net4 vss 87.3011e-18
c2966 n581__r_out vss 197.806e-18
c2967 n585__r_out vss 80.9816e-18
c2968 n477__i18__net5 vss 61.12e-21
c2969 n14__i14__i17__i2__net5 vss 143.359e-18
c2970 n14__i14__i17__i3__net5 vss 143.078e-18
c2971 n354__vddio vss 129.729e-18
c2972 n355__vddio vss 122.73e-18
c2973 n358__vddio vss 109.373e-18
c2974 n359__vddio vss 82.4675e-18
c2975 n9__i14__i13__net4 vss 76.7283e-18
c2976 n9__i14__i16__net4 vss 76.4897e-18
c2977 n9__i14__i10__net4 vss 74.3248e-18
c2978 n9__i14__i9__net4 vss 73.4915e-18
c2979 n12__i14__i13__net4 vss 113.903e-18
c2980 n12__i14__i16__net4 vss 113.815e-18
c2981 n12__i14__i10__net4 vss 113.978e-18
c2982 n12__i14__i9__net4 vss 113.721e-18
c2983 n10__i14__i17__net6 vss 466.814e-18
c2984 n11__i14__i17__net6 vss 454.271e-18
c2985 n475__i18__net5 vss 61.12e-21
c2986 n568__r_out vss 131.6e-18
c2987 n572__r_out vss 79.0526e-18
c2988 n14__i14__i13__net5 vss 138.422e-18
c2989 n14__i14__i16__net5 vss 138.703e-18
c2990 n14__i14__i10__net5 vss 137.982e-18
c2991 n14__i14__i9__net5 vss 139.264e-18
c2992 n473__i18__net5 vss 61.12e-21
c2993 n17__i14__net4 vss 75.867e-18
c2994 n18__i14__net4 vss 71.9878e-18
c2995 n19__i14__net4 vss 72.4663e-18
c2996 n20__i14__net4 vss 69.8719e-18
c2997 n7__i14__i17__i2__net4 vss 150.613e-18
c2998 n7__i14__i17__i3__net4 vss 156.678e-18
c2999 n345__vddio vss 135.666e-18
c3000 n348__vddio vss 115.33e-18
c3001 n349__vddio vss 113.768e-18
c3002 n352__vddio vss 86.1419e-18
c3003 n468__i18__net5 vss 61.12e-21
c3004 n11__i14__i17__i2__net5 vss 116.574e-18
c3005 n11__i14__i17__i3__net5 vss 115.952e-18
c3006 n1__vdd vss 117.467e-18
c3007 n4__vdd vss 159.493e-18
c3008 n5__vdd vss 240.936e-18
c3009 n555__r_out vss 131.608e-18
c3010 n559__r_out vss 74.4276e-18
c3011 n7__i14__i13__net4 vss 173.583e-18
c3012 n7__i14__i16__net4 vss 173.675e-18
c3013 n7__i14__i10__net4 vss 173.759e-18
c3014 n7__i14__i9__net4 vss 173.458e-18
c3015 n21__ck vss 199.94e-18
c3016 n11__i14__i17__net3 vss 195.01e-18
c3017 n20__i14__i17__net1 vss 189.737e-18
c3018 n12__i14__i17__net7 vss 198.789e-18
c3019 n467__i18__net5 vss 61.12e-21
c3020 n338__vddio vss 127.669e-18
c3021 n339__vddio vss 121.868e-18
c3022 n342__vddio vss 108.044e-18
c3023 n343__vddio vss 80.4072e-18
c3024 n11__i14__i13__net5 vss 119.479e-18
c3025 n11__i14__i16__net5 vss 120.023e-18
c3026 n11__i14__i10__net5 vss 119.668e-18
c3027 n11__i14__i9__net5 vss 120.112e-18
c3028 n461__i18__net5 vss 61.12e-21
c3029 n53__i14__net10 vss 195.585e-18
c3030 n45__i14__net9 vss 170.248e-18
c3031 n46__i14__net9 vss 170.129e-18
c3032 n54__i14__net10 vss 195.521e-18
c3033 n55__i14__net10 vss 199.248e-18
c3034 n47__i14__net9 vss 170.149e-18
c3035 n48__i14__net9 vss 170.238e-18
c3036 n56__i14__net10 vss 195.655e-18
c3037 n542__r_out vss 203.417e-18
c3038 n546__r_out vss 73.0572e-18
c3039 n5__i14__i17__i2__net2 vss 205.545e-18
c3040 n5__i14__i17__i3__net2 vss 213.093e-18
c3041 n456__i18__net5 vss 61.12e-21
c3042 n330__vddio vss 131.014e-18
c3043 n331__vddio vss 124.577e-18
c3044 n334__vddio vss 110.302e-18
c3045 n335__vddio vss 83.7851e-18
c3046 n16__i14__i17__i2__net1 vss 113.832e-18
c3047 n16__i14__i17__i3__net1 vss 113.769e-18
c3048 n5__i14__i13__net2 vss 209.427e-18
c3049 n5__i14__i16__net2 vss 209.43e-18
c3050 n5__i14__i10__net2 vss 209.415e-18
c3051 n5__i14__i9__net2 vss 209.422e-18
c3052 n449__i18__net5 vss 61.12e-21
c3053 n19__reset vss 285.029e-18
c3054 n14__i14__i17__i2__net1 vss 256.58e-18
c3055 n14__i14__i17__i3__net1 vss 256.955e-18
c3056 n529__r_out vss 130.842e-18
c3057 n533__r_out vss 78.5259e-18
c3058 n10__i14__i17__net3 vss 329.126e-18
c3059 n19__i14__i17__net1 vss 327.864e-18
c3060 n446__i18__net5 vss 61.12e-21
c3061 n16__i14__i13__net1 vss 113.783e-18
c3062 n16__i14__i16__net1 vss 113.983e-18
c3063 n16__i14__i10__net1 vss 113.585e-18
c3064 n16__i14__i9__net1 vss 113.902e-18
c3065 n15__ck vss 287.647e-18
c3066 n16__ck vss 250.095e-18
c3067 n10__i14__i17__net7 vss 188.775e-18
c3068 n11__i14__i17__net7 vss 287.989e-18
c3069 n10__i14__net3 vss 523.175e-18
c3070 n11__i14__net3 vss 513.987e-18
c3071 n322__vddio vss 131.013e-18
c3072 n323__vddio vss 123.674e-18
c3073 n326__vddio vss 110.302e-18
c3074 n327__vddio vss 83.7851e-18
c3075 n14__i14__i13__net1 vss 257.362e-18
c3076 n14__i14__i16__net1 vss 256.839e-18
c3077 n14__i14__i10__net1 vss 257.226e-18
c3078 n14__i14__i9__net1 vss 256.934e-18
c3079 n9__i14__i17__net3 vss 271.628e-18
c3080 n18__i14__i17__net1 vss 259.1e-18
c3081 n438__i18__net5 vss 61.12e-21
c3082 n41__i14__net9 vss 325.856e-18
c3083 n42__i14__net9 vss 325.236e-18
c3084 n43__i14__net9 vss 325.642e-18
c3085 n44__i14__net9 vss 325.028e-18
c3086 n514__r_out vss 205.05e-18
c3087 n515__r_out vss 78.7721e-18
c3088 n49__i14__net10 vss 302.509e-18
c3089 n37__i14__net10 vss 255.107e-18
c3090 n50__i14__net10 vss 285.511e-18
c3091 n51__i14__net10 vss 285.914e-18
c3092 n41__i14__net10 vss 237.607e-18
c3093 n52__i14__net10 vss 284.808e-18
c3094 n4__i14__i17__i2__net2 vss 240.666e-18
c3095 n4__i14__i17__i3__net2 vss 243.544e-18
c3096 n434__i18__net5 vss 61.12e-21
c3097 n21__i14__net9 vss 290.499e-18
c3098 n25__i14__net9 vss 269.489e-18
c3099 n314__vddio vss 127.671e-18
c3100 n315__vddio vss 120.899e-18
c3101 n318__vddio vss 108.044e-18
c3102 n319__vddio vss 80.4072e-18
c3103 n11__i14__i17__i2__net1 vss 247.036e-18
c3104 n11__i14__i17__i3__net1 vss 245.087e-18
c3105 n431__i18__net5 vss 61.12e-21
c3106 n13__ck vss 158.143e-18
c3107 n7__i14__i17__net7 vss 88.3111e-18
c3108 n4__i14__i13__net2 vss 242.867e-18
c3109 n4__i14__i16__net2 vss 242.932e-18
c3110 n4__i14__i10__net2 vss 242.886e-18
c3111 n4__i14__i9__net2 vss 242.908e-18
c3112 n8__i14__i17__net3 vss 243.196e-18
c3113 n10__i14__i17__net1 vss 162.671e-18
c3114 n501__r_out vss 64.6114e-18
c3115 n502__r_out vss 78.2152e-18
c3116 n6__i14__i17__net1 vss 141.603e-18
c3117 n2__i14__i17__net8 vss 129.644e-18
c3118 n11__i14__i13__net1 vss 240.652e-18
c3119 n11__i14__i16__net1 vss 240.13e-18
c3120 n11__i14__i10__net1 vss 240.484e-18
c3121 n11__i14__i9__net1 vss 240.557e-18
c3122 n426__i18__net5 vss 61.12e-21
c3123 n6__i14__i17__net3 vss 137.576e-18
c3124 n6__i14__i17__net6 vss 112.591e-18
c3125 n18__i14__net10 vss 145.871e-18
c3126 n22__i14__net10 vss 145.065e-18
c3127 n24__i14__net10 vss 145.777e-18
c3128 n28__i14__net10 vss 145.516e-18
c3129 n306__vddio vss 127.671e-18
c3130 n307__vddio vss 121.142e-18
c3131 n310__vddio vss 108.044e-18
c3132 n311__vddio vss 80.4072e-18
c3133 n17__i14__net9 vss 262.6e-18
c3134 n18__i14__net9 vss 256.275e-18
c3135 n19__i14__net9 vss 257.143e-18
c3136 n20__i14__net9 vss 257.113e-18
c3137 n8__ck vss 48.9541e-18
c3138 n418__i18__net5 vss 61.12e-21
c3139 n2__x3 vss 80.9545e-18
c3140 n2__x2 vss 79.7459e-18
c3141 n2__x1 vss 176.336e-18
c3142 n2__x0 vss 176.3e-18
c3143 n487__r_out vss 125.772e-18
c3144 n490__r_out vss 84.8543e-18
c3145 n416__i18__net5 vss 61.12e-21
c3146 n298__vddio vss 129.727e-18
c3147 n299__vddio vss 122.82e-18
c3148 n302__vddio vss 109.373e-18
c3149 n303__vddio vss 82.4675e-18
c3150 n411__i18__net5 vss 61.12e-21
c3151 n474__r_out vss 199.397e-18
c3152 n477__r_out vss 85.0746e-18
c3153 n403__i18__net5 vss 61.12e-21
c3154 n290__vddio vss 129.729e-18
c3155 n291__vddio vss 122.73e-18
c3156 n294__vddio vss 109.373e-18
c3157 n295__vddio vss 82.4675e-18
c3158 n402__i18__net5 vss 61.12e-21
c3159 n464__r_out vss 58.5197e-18
c3160 n468__r_out vss 85.7165e-18
c3161 n393__i18__net5 vss 61.12e-21
c3162 n282__vddio vss 127.671e-18
c3163 n283__vddio vss 121.052e-18
c3164 n286__vddio vss 108.044e-18
c3165 n287__vddio vss 80.4072e-18
c3166 n388__i18__net5 vss 61.12e-21
c3167 n448__r_out vss 59.85e-18
c3168 n452__r_out vss 85.3776e-18
c3169 n383__i18__net5 vss 61.12e-21
c3170 n274__vddio vss 127.671e-18
c3171 n275__vddio vss 121.868e-18
c3172 n278__vddio vss 108.044e-18
c3173 n279__vddio vss 80.4072e-18
c3174 n381__i18__net5 vss 61.12e-21
c3175 n432__r_out vss 58.7858e-18
c3176 n435__r_out vss 83.9817e-18
c3177 n373__i18__net5 vss 61.12e-21
c3178 n266__vddio vss 131.014e-18
c3179 n267__vddio vss 124.577e-18
c3180 n270__vddio vss 110.302e-18
c3181 n271__vddio vss 83.7851e-18
c3182 n371__i18__net5 vss 61.12e-21
c3183 n420__r_out vss 59.0518e-18
c3184 n424__r_out vss 85.2875e-18
c3185 n363__i18__net5 vss 61.12e-21
c3186 n258__vddio vss 131.012e-18
c3187 n259__vddio vss 123.674e-18
c3188 n262__vddio vss 110.302e-18
c3189 n263__vddio vss 83.7851e-18
c3190 n358__i18__net5 vss 61.12e-21
c3191 n407__r_out vss 59.85e-18
c3192 n411__r_out vss 85.5795e-18
c3193 n353__i18__net5 vss 61.12e-21
c3194 n250__vddio vss 127.671e-18
c3195 n251__vddio vss 120.914e-18
c3196 n254__vddio vss 108.044e-18
c3197 n255__vddio vss 80.4072e-18
c3198 n351__i18__net5 vss 61.12e-21
c3199 n391__r_out vss 58.7858e-18
c3200 n394__r_out vss 84.7417e-18
c3201 n343__i18__net5 vss 61.12e-21
c3202 n242__vddio vss 129.729e-18
c3203 n243__vddio vss 122.82e-18
c3204 n246__vddio vss 109.373e-18
c3205 n247__vddio vss 82.4675e-18
c3206 n341__i18__net5 vss 61.12e-21
c3207 n378__r_out vss 199.186e-18
c3208 n381__r_out vss 85.075e-18
c3209 n333__i18__net5 vss 61.12e-21
c3210 n234__vddio vss 129.729e-18
c3211 n235__vddio vss 122.73e-18
c3212 n238__vddio vss 109.373e-18
c3213 n239__vddio vss 82.4675e-18
c3214 n331__i18__net5 vss 61.12e-21
c3215 n365__r_out vss 58.7858e-18
c3216 n368__r_out vss 86.0029e-18
c3217 n323__i18__net5 vss 61.12e-21
c3218 n226__vddio vss 127.671e-18
c3219 n227__vddio vss 121.052e-18
c3220 n230__vddio vss 108.044e-18
c3221 n231__vddio vss 80.4072e-18
c3222 n318__i18__net5 vss 61.12e-21
c3223 n352__r_out vss 198.935e-18
c3224 n355__r_out vss 85.1891e-18
c3225 n316__i18__net5 vss 61.12e-21
c3226 n218__vddio vss 127.669e-18
c3227 n219__vddio vss 121.868e-18
c3228 n222__vddio vss 108.044e-18
c3229 n223__vddio vss 80.4072e-18
c3230 n308__i18__net5 vss 61.12e-21
c3231 n342__r_out vss 198.781e-18
c3232 n346__r_out vss 83.9519e-18
c3233 n306__i18__net5 vss 61.12e-21
c3234 n210__vddio vss 131.014e-18
c3235 n211__vddio vss 124.735e-18
c3236 n214__vddio vss 110.302e-18
c3237 n215__vddio vss 83.7851e-18
c3238 n301__i18__net5 vss 61.12e-21
c3239 n326__r_out vss 58.7858e-18
c3240 n329__r_out vss 85.1878e-18
c3241 n296__i18__net5 vss 61.12e-21
c3242 n202__vddio vss 131.014e-18
c3243 n203__vddio vss 123.674e-18
c3244 n206__vddio vss 110.302e-18
c3245 n207__vddio vss 83.7851e-18
c3246 n291__i18__net5 vss 61.12e-21
c3247 n313__r_out vss 59.85e-18
c3248 n316__r_out vss 85.595e-18
c3249 n286__i18__net5 vss 61.12e-21
c3250 n194__vddio vss 127.671e-18
c3251 n195__vddio vss 120.899e-18
c3252 n198__vddio vss 108.044e-18
c3253 n199__vddio vss 80.4072e-18
c3254 n281__i18__net5 vss 61.12e-21
c3255 n300__r_out vss 58.7858e-18
c3256 n303__r_out vss 85.0284e-18
c3257 n273__i18__net5 vss 61.12e-21
c3258 n186__vddio vss 127.671e-18
c3259 n187__vddio vss 121.142e-18
c3260 n190__vddio vss 108.044e-18
c3261 n191__vddio vss 80.4072e-18
c3262 n271__i18__net5 vss 61.12e-21
c3263 n287__r_out vss 59.0518e-18
c3264 n290__r_out vss 84.9217e-18
c3265 n263__i18__net5 vss 61.12e-21
c3266 n178__vddio vss 129.727e-18
c3267 n179__vddio vss 122.82e-18
c3268 n182__vddio vss 109.373e-18
c3269 n183__vddio vss 82.4675e-18
c3270 n261__i18__net5 vss 61.12e-21
c3271 n277__r_out vss 59.85e-18
c3272 n281__r_out vss 85.1453e-18
c3273 n256__i18__net5 vss 61.12e-21
c3274 n170__vddio vss 129.729e-18
c3275 n171__vddio vss 122.73e-18
c3276 n174__vddio vss 109.373e-18
c3277 n175__vddio vss 82.4675e-18
c3278 n248__i18__net5 vss 61.12e-21
c3279 n261__r_out vss 58.7858e-18
c3280 n264__r_out vss 85.6422e-18
c3281 n243__i18__net5 vss 61.12e-21
c3282 n162__vddio vss 127.671e-18
c3283 n163__vddio vss 121.052e-18
c3284 n166__vddio vss 108.044e-18
c3285 n167__vddio vss 80.4072e-18
c3286 n238__i18__net5 vss 61.12e-21
c3287 n248__r_out vss 59.85e-18
c3288 n251__r_out vss 85.3702e-18
c3289 n233__i18__net5 vss 61.12e-21
c3290 n154__vddio vss 127.671e-18
c3291 n155__vddio vss 121.868e-18
c3292 n158__vddio vss 108.044e-18
c3293 n159__vddio vss 80.4072e-18
c3294 n231__i18__net5 vss 61.12e-21
c3295 n235__r_out vss 58.7907e-18
c3296 n238__r_out vss 82.3621e-18
c3297 n226__i18__net5 vss 122.24e-21
c3298 n146__vddio vss 131.214e-18
c3299 n147__vddio vss 125.11e-18
c3300 n150__vddio vss 110.43e-18
c3301 n151__vddio vss 83.7851e-18
c3302 n221__i18__net5 vss 122.24e-21
c3303 n222__r_out vss 59.0567e-18
c3304 n225__r_out vss 82.8563e-18
c3305 n213__i18__net5 vss 122.24e-21
c3306 n138__vddio vss 131.214e-18
c3307 n139__vddio vss 124.197e-18
c3308 n142__vddio vss 110.43e-18
c3309 n143__vddio vss 83.7851e-18
c3310 n211__i18__net5 vss 122.24e-21
c3311 n212__r_out vss 59.8549e-18
c3312 n216__r_out vss 83.1529e-18
c3313 n206__i18__net5 vss 122.24e-21
c3314 n130__vddio vss 127.818e-18
c3315 n131__vddio vss 121.343e-18
c3316 n134__vddio vss 108.172e-18
c3317 n135__vddio vss 80.4072e-18
c3318 n198__i18__net5 vss 122.24e-21
c3319 n196__r_out vss 58.7907e-18
c3320 n199__r_out vss 82.9261e-18
c3321 n196__i18__net5 vss 985.066e-21
c3322 n122__vddio vss 129.108e-18
c3323 n123__vddio vss 122.249e-18
c3324 n126__vddio vss 108.835e-18
c3325 n127__vddio vss 81.6979e-18
c3326 n191__i18__net5 vss 122.24e-21
c3327 n183__r_out vss 196.449e-18
c3328 n186__r_out vss 82.6119e-18
c3329 n183__i18__net5 vss 5.16372e-18
c3330 n114__vddio vss 129.108e-18
c3331 n115__vddio vss 122.062e-18
c3332 n118__vddio vss 108.835e-18
c3333 n119__vddio vss 81.6979e-18
c3334 n178__i18__net5 vss 122.24e-21
c3335 n170__r_out vss 58.7907e-18
c3336 n173__r_out vss 83.3845e-18
c3337 n176__i18__net5 vss 349.913e-21
c3338 n106__vddio vss 130.836e-18
c3339 n107__vddio vss 123.863e-18
c3340 n110__vddio vss 110.163e-18
c3341 n111__vddio vss 83.408e-18
c3342 n168__i18__net5 vss 204.81e-21
c3343 n157__r_out vss 199.464e-18
c3344 n160__r_out vss 82.2281e-18
c3345 n163__i18__net5 vss 122.24e-21
c3346 n98__vddio vss 130.836e-18
c3347 n99__vddio vss 124.801e-18
c3348 n102__vddio vss 110.163e-18
c3349 n103__vddio vss 83.408e-18
c3350 n158__i18__net5 vss 122.24e-21
c3351 n147__r_out vss 199.261e-18
c3352 n151__r_out vss 81.5436e-18
c3353 n156__i18__net5 vss 122.24e-21
c3354 n90__vddio vss 129.88e-18
c3355 n91__vddio vss 124.026e-18
c3356 n94__vddio vss 109.501e-18
c3357 n95__vddio vss 82.4675e-18
c3358 n151__i18__net5 vss 122.24e-21
c3359 n134__r_out vss 58.7907e-18
c3360 n138__r_out vss 82.8416e-18
c3361 n146__i18__net5 vss 122.24e-21
c3362 n82__vddio vss 129.204e-18
c3363 n83__vddio vss 122.512e-18
c3364 n86__vddio vss 109.157e-18
c3365 n87__vddio vss 82.4675e-18
c3366 n141__i18__net5 vss 61.12e-21
c3367 n118__r_out vss 59.85e-18
c3368 n121__r_out vss 85.7623e-18
c3369 n133__i18__net5 vss 61.12e-21
c3370 n74__vddio vss 127.671e-18
c3371 n75__vddio vss 121.052e-18
c3372 n78__vddio vss 108.044e-18
c3373 n79__vddio vss 80.4072e-18
c3374 n128__i18__net5 vss 61.12e-21
c3375 n105__r_out vss 58.7858e-18
c3376 n108__r_out vss 84.9114e-18
c3377 n126__i18__net5 vss 61.12e-21
c3378 n66__vddio vss 126.946e-18
c3379 n67__vddio vss 120.583e-18
c3380 n70__vddio vss 107.485e-18
c3381 n71__vddio vss 80.3408e-18
c3382 n119__i18__net5 vss 61.12e-21
c3383 n92__r_out vss 59.0518e-18
c3384 n95__r_out vss 82.3896e-18
c3385 n113__i18__net5 vss 61.12e-21
c3386 n58__vddio vss 128.744e-18
c3387 n59__vddio vss 121.73e-18
c3388 n62__vddio vss 108.623e-18
c3389 n63__vddio vss 81.6878e-18
c3390 n109__i18__net5 vss 61.12e-21
c3391 n82__r_out vss 59.85e-18
c3392 n86__r_out vss 82.7715e-18
c3393 n106__i18__net5 vss 61.12e-21
c3394 n50__vddio vss 128.744e-18
c3395 n51__vddio vss 121.485e-18
c3396 n54__vddio vss 108.623e-18
c3397 n55__vddio vss 81.6878e-18
c3398 n98__i18__net5 vss 61.12e-21
c3399 n66__r_out vss 58.7858e-18
c3400 n69__r_out vss 83.1156e-18
c3401 n93__i18__net5 vss 61.12e-21
c3402 n42__vddio vss 130.449e-18
c3403 n43__vddio vss 123.242e-18
c3404 n46__vddio vss 109.943e-18
c3405 n47__vddio vss 83.3979e-18
c3406 n88__i18__net5 vss 61.12e-21
c3407 n53__r_out vss 199.373e-18
c3408 n56__r_out vss 82.4599e-18
c3409 n83__i18__net5 vss 61.12e-21
c3410 n34__vddio vss 130.449e-18
c3411 n35__vddio vss 124.169e-18
c3412 n38__vddio vss 109.943e-18
c3413 n39__vddio vss 83.3979e-18
c3414 n81__i18__net5 vss 61.12e-21
c3415 n40__r_out vss 58.7858e-18
c3416 n43__r_out vss 81.7292e-18
c3417 n76__i18__net5 vss 61.12e-21
c3418 n26__vddio vss 129.511e-18
c3419 n27__vddio vss 123.428e-18
c3420 n30__vddio vss 109.282e-18
c3421 n31__vddio vss 82.4574e-18
c3422 n71__i18__net5 vss 61.12e-21
c3423 n27__r_out vss 199.469e-18
c3424 n30__r_out vss 82.9643e-18
c3425 n66__i18__net5 vss 61.12e-21
c3426 n18__vddio vss 129.511e-18
c3427 n19__vddio vss 122.636e-18
c3428 n22__vddio vss 109.282e-18
c3429 n23__vddio vss 82.4574e-18
c3430 n58__i18__net5 vss 61.12e-21
c3431 n17__r_out vss 199.099e-18
c3432 n21__r_out vss 83.5087e-18
c3433 n56__i18__net5 vss 404.265e-21
c3434 n10__vddio vss 127.818e-18
c3435 n11__vddio vss 121.292e-18
c3436 n14__vddio vss 108.266e-18
c3437 n15__vddio vss 80.6068e-18
c3438 n48__i18__net5 vss 61.12e-21
c3439 n1__r_out vss 58.7837e-18
c3440 n4__r_out vss 85.1035e-18
c3441 n46__i18__net5 vss 7.18615e-18
c3442 n2__vddio vss 71.927e-18
c3443 n3__vddio vss 68.3216e-18
c3444 n6__vddio vss 60.6355e-18
c3445 n7__vddio vss 51.7365e-18
c3446 n686__vddio vss 27.7472e-15
c3447 n683__vddio vss 133.561e-18
c3448 n678__vddio vss 127.285e-18
c3449 n9__i18__net1 vss 135.968e-18
c3450 n8__r0_buff vss 35.6963e-18
c3451 n8__r2_buff vss 43.2132e-18
c3452 n8__r1_buff vss 43.2132e-18
c3453 n133__vdd vss 62.5539e-18
c3454 n291__vdd vss 64.1374e-18
c3455 n349__vdd vss 64.1417e-18
c3456 n7__serial_out_b_high_buff vss 126.664e-18
c3457 n14__r0_buff vss 57.3722e-18
c3458 n14__r2_buff vss 57.423e-18
c3459 n14__r1_buff vss 57.1623e-18
c3460 n685__vddio vss 72.3027e-18
c3461 n211__vdd vss 55.3399e-18
c3462 n351__vdd vss 57.2577e-18
c3463 n350__vdd vss 57.2577e-18
c3464 n7__i18__net1 vss 117.831e-18
c3465 n13__r1_buff vss 48.5352e-21
c3466 n6__serial_out_b_high_buff vss 106.294e-18
c3467 n134__vdd vss 2.52778e-15
c3468 n293__vdd vss 3.08678e-15
c3469 n11__r0_buff vss 31.7017e-18
c3470 n15__r2_buff vss 30.9089e-18
c3471 n11__r1_buff vss 32.5376e-18
c3472 n12__net7 vss 29.862e-18
c3473 n13__net6 vss 29.4732e-18
c3474 n12__net8 vss 29.8977e-18
c3475 n132__vdd vss 28.512e-18
c3476 n11__i12__bcore_bar vss 34.0122e-18
c3477 n13__net7 vss 45.9376e-18
c3478 n12__net6 vss 45.9783e-18
c3479 n13__net8 vss 45.4917e-18
c3480 n130__vdd vss 36.8889e-18
c3481 n682__vddio vss 112.113e-18
c3482 n212__vdd vss 40.4343e-18
c3483 n353__vdd vss 47.6557e-18
c3484 n352__vdd vss 47.2921e-18
c3485 n14__i12__bcore_bar vss 52.313e-18
c3486 n15__i18__net2 vss 283.475e-18
c3487 n681__vddio vss 168.908e-18
c3488 n676__vddio vss 52.3589e-18
c3489 n659__vddio vss 283.667e-18
c3490 n5__i12__bio vss 41.6288e-18
c3491 n3__i1__q vss 76.744e-18
c3492 n56__i18__net3 vss 498.459e-18
c3493 n213__vdd vss 90.2167e-18
c3494 n355__vdd vss 89.8531e-18
c3495 n354__vdd vss 90.3114e-18
c3496 n23__serial_out vss 56.3843e-18
c3497 n14__net4 vss 60.1325e-18
c3498 n13__net3 vss 61.0279e-18
c3499 n664__vddio vss 486.092e-18
c3500 n214__vdd vss 62.5355e-18
c3501 n357__vdd vss 64.3982e-18
c3502 n356__vdd vss 65.8887e-18
c3503 n677__vddio vss 53.7218e-18
c3504 n58__i18__net3 vss 495.819e-18
c3505 n215__vdd vss 56.4903e-18
c3506 n359__vdd vss 58.1182e-18
c3507 n358__vdd vss 58.3752e-18
c3508 n6__serial_out_b_high vss 25.8079e-18
c3509 n10__i2__net77 vss 45.2955e-18
c3510 n10__i1__net77 vss 45.6196e-18
c3511 n10__i0__net77 vss 45.4371e-18
c3512 n662__vddio vss 290.249e-18
c3513 n216__vdd vss 91.4789e-18
c3514 n361__vdd vss 93.1705e-18
c3515 n360__vdd vss 93.923e-18
c3516 n15__i2__net76 vss 16.8525e-21
c3517 n15__i1__net76 vss 16.8525e-21
c3518 n15__i0__net76 vss 16.8525e-21
c3519 n217__vdd vss 26.4412e-18
c3520 n363__vdd vss 27.5141e-18
c3521 n362__vdd vss 26.1499e-18
c3522 n636__vddio vss 403.122e-18
c3523 n218__vdd vss 51.6434e-18
c3524 n365__vdd vss 52.134e-18
c3525 n364__vdd vss 49.8557e-18
c3526 n10__r1 vss 39.0164e-18
c3527 n26__i13__net18 vss 82.0488e-18
c3528 n200__i18__net4 vss 636.3e-18
c3529 n9__i2__net76 vss 37.9914e-18
c3530 n9__i1__net76 vss 39.9866e-18
c3531 n9__i0__net76 vss 38.4885e-18
c3532 n643__vddio vss 686.777e-18
c3533 n13__i2__net76 vss 84.0604e-18
c3534 n12__i1__net76 vss 93.5967e-18
c3535 n13__i0__net76 vss 94.5181e-18
c3536 n6__i2__net75 vss 81.8608e-18
c3537 n11__i1__net75 vss 87.8736e-18
c3538 n6__i0__net75 vss 88.9805e-18
c3539 n189__i18__net4 vss 640.105e-18
c3540 n5__i13__i20__i4__net2 vss 112.936e-18
c3541 n219__vdd vss 93.5695e-18
c3542 n367__vdd vss 91.8793e-18
c3543 n366__vdd vss 95.4638e-18
c3544 n68__vdd vss 72.9741e-18
c3545 n11__i2__net75 vss 48.8317e-18
c3546 n9__i1__net75 vss 48.5471e-18
c3547 n11__i0__net75 vss 48.6937e-18
c3548 n646__vddio vss 690.564e-18
c3549 n220__vdd vss 98.2441e-18
c3550 n369__vdd vss 97.602e-18
c3551 n368__vdd vss 97.9655e-18
c3552 n9__i13__net23 vss 70.2609e-18
c3553 n183__i18__net4 vss 640.105e-18
c3554 n70__vdd vss 70.9344e-18
c3555 n69__vdd vss 63.2609e-18
c3556 n653__vddio vss 690.375e-18
c3557 n10__i13__i20__net1 vss 75.1484e-18
c3558 n7__i13__net3 vss 94.6481e-18
c3559 n71__vdd vss 58.1564e-18
c3560 n167__i18__net4 vss 640.148e-18
c3561 n72__vdd vss 80.8469e-18
c3562 n221__vdd vss 94.8777e-18
c3563 n371__vdd vss 95.0359e-18
c3564 n370__vdd vss 93.5119e-18
c3565 n656__vddio vss 749.205e-18
c3566 n9__i2__net74 vss 39.2111e-18
c3567 n9__i1__net74 vss 42.7627e-18
c3568 n9__i0__net74 vss 39.588e-18
c3569 n156__i18__net4 vss 650.679e-18
c3570 n13__i2__net74 vss 86.0367e-18
c3571 n12__i1__net74 vss 98.6319e-18
c3572 n13__i0__net74 vss 97.1819e-18
c3573 n5__i1__net73 vss 80.3804e-18
c3574 n650__vddio vss 425.383e-18
c3575 n16__i13__net18 vss 39.2494e-18
c3576 n5__r0 vss 37.1943e-18
c3577 n13__i18__net2 vss 219.566e-18
c3578 n672__vddio vss 205.738e-18
c3579 n9__i12__bio vss 51.9544e-18
c3580 n3__i2__q vss 46.4112e-18
c3581 n3__i0__q vss 43.4022e-18
c3582 n51__i18__net3 vss 375.375e-18
c3583 n21__serial_out vss 55.3102e-18
c3584 n15__net4 vss 54.1916e-18
c3585 n11__net3 vss 53.9671e-18
c3586 n3__i12__bio vss 42.997e-18
c3587 n60__i18__net3 vss 373.385e-18
c3588 n8__i2__net77 vss 65.9037e-18
c3589 n8__i1__net77 vss 65.2606e-18
c3590 n8__i0__net77 vss 63.8647e-18
c3591 n8__serial_out_b_high vss 124.56e-18
c3592 n32__vdd vss 3.53512e-15
c3593 n9__r1 vss 53.8915e-18
c3594 n10__serial_out_b_high vss 118.543e-18
c3595 n196__i18__net4 vss 464.651e-18
c3596 n8__i2__net76 vss 37.8293e-18
c3597 n8__i1__net76 vss 36.1873e-18
c3598 n8__i0__net76 vss 37.7128e-18
c3599 n5__r1 vss 103.947e-18
c3600 n12__i2__net76 vss 58.8165e-18
c3601 n13__i1__net76 vss 57.7253e-18
c3602 n12__i0__net76 vss 55.8034e-18
c3603 n16__i13__net7 vss 90.0591e-18
c3604 n10__i2__net75 vss 36.0303e-18
c3605 n6__i1__net75 vss 36.1071e-18
c3606 n10__i0__net75 vss 34.2841e-18
c3607 n185__i18__net4 vss 464.979e-18
c3608 n3__i13__i20__i4__net2 vss 21.9217e-18
c3609 n9__i2__net75 vss 64.4665e-18
c3610 n12__i1__net75 vss 63.4077e-18
c3611 n9__i0__net75 vss 59.1416e-18
c3612 n7__i13__net23 vss 38.8968e-18
c3613 n3__r2 vss 30.9789e-18
c3614 n180__i18__net4 vss 464.81e-18
c3615 n14__i2__net74 vss 61.8044e-18
c3616 n14__i1__net74 vss 62.51e-18
c3617 n14__i0__net74 vss 65.5511e-18
c3618 n8__i13__i20__net1 vss 69.2111e-18
c3619 n9__i13__net3 vss 58.5752e-18
c3620 n163__i18__net4 vss 463.764e-18
c3621 n8__i2__net74 vss 36.7269e-18
c3622 n8__i1__net74 vss 36.7913e-18
c3623 n8__i0__net74 vss 36.3531e-18
c3624 n152__i18__net4 vss 472.269e-18
c3625 n12__i2__net74 vss 59.4356e-18
c3626 n13__i1__net74 vss 58.9059e-18
c3627 n12__i0__net74 vss 56.1102e-18
c3628 n5__i2__net73 vss 25.5479e-18
c3629 n5__i0__net73 vss 26.301e-18
c3630 n15__i13__net18 vss 54.621e-18
c3631 n8__r0 vss 53.0539e-18
c3632 n22__i13__net1 vss 82.5325e-18
c3633 n26__i13__net2 vss 81.8053e-18
c3634 n6__i2__net73 vss 75.344e-18
c3635 n4__i1__net73 vss 81.3878e-18
c3636 n6__i0__net73 vss 78.9844e-18
c3637 n5__i13__i19__i4__net2 vss 112.804e-18
c3638 n3__i13__i18__i4__net2 vss 112.427e-18
c3639 n222__vdd vss 86.7177e-18
c3640 n373__vdd vss 1.02474e-18
c3641 n372__vdd vss 1.04156e-18
c3642 n535__vddio vss 282.599e-18
c3643 n74__vdd vss 74.3623e-18
c3644 n73__vdd vss 74.3818e-18
c3645 n689__i18__net5 vss 883.924e-18
c3646 n8__i13__net17 vss 71.0467e-18
c3647 n12__i13__net7 vss 71.089e-18
c3648 n76__vdd vss 67.3869e-18
c3649 n75__vdd vss 67.8654e-18
c3650 n560__vddio vss 464.594e-18
c3651 n3__r0_buff vss 52.892e-18
c3652 n3__r1_buff vss 51.3416e-18
c3653 n3__r2_buff vss 51.6693e-18
c3654 n10__i13__i19__net1 vss 77.6728e-18
c3655 n10__i13__i18__net1 vss 77.192e-18
c3656 n5__i2__net1 vss 273.45e-18
c3657 n5__i1__net1 vss 272.292e-18
c3658 n5__i0__net1 vss 271.444e-18
c3659 n681__i18__net5 vss 825.624e-18
c3660 n78__vdd vss 57.543e-18
c3661 n77__vdd vss 57.4285e-18
c3662 n4__net4 vss 68.7037e-18
c3663 n4__net3 vss 67.6138e-18
c3664 n564__vddio vss 462.79e-18
c3665 n9__i2__net79 vss 51.7163e-18
c3666 n9__i1__net79 vss 53.074e-18
c3667 n9__i0__net79 vss 53.3753e-18
c3668 n223__vdd vss 40.8137e-18
c3669 n375__vdd vss 46.0714e-18
c3670 n374__vdd vss 47.0316e-18
c3671 n663__i18__net5 vss 832.129e-18
c3672 n224__vdd vss 46.799e-18
c3673 n568__vddio vss 462.874e-18
c3674 n29__shift vss 51.052e-18
c3675 n14__i13__net12 vss 47.25e-18
c3676 n15__i13__net2 vss 46.0896e-18
c3677 n225__vdd vss 87.7777e-18
c3678 n650__i18__net5 vss 830.415e-18
c3679 n28__i13__a2 vss 82.4554e-18
c3680 n28__i13__a0 vss 82.4576e-18
c3681 n25__shift vss 49.6329e-18
c3682 n15__reset_buff vss 54.4002e-18
c3683 n572__vddio vss 462.915e-18
c3684 n376__vdd vss 104.548e-18
c3685 n226__vdd vss 68.1747e-18
c3686 n12__reset_buff vss 69.5474e-18
c3687 n642__i18__net5 vss 830.94e-18
c3688 n377__vdd vss 76.8235e-18
c3689 n5__i13__i17__i4__net2 vss 114.367e-18
c3690 n3__i13__i16__i4__net2 vss 113.972e-18
c3691 n7__i9__net1 vss 79.1237e-18
c3692 n11__i13__net18 vss 106.491e-18
c3693 n16__i13__net11 vss 89.7513e-18
c3694 n20__i13__net12 vss 89.345e-18
c3695 n4__i2__net73 vss 52.9943e-18
c3696 n6__i1__net73 vss 52.8177e-18
c3697 n4__i0__net73 vss 49.2948e-18
c3698 n3__i13__i19__i4__net2 vss 22.0092e-18
c3699 n5__i13__i18__i4__net2 vss 285.033e-21
c3700 n684__i18__net5 vss 616.736e-18
c3701 n6__i13__net17 vss 40.7179e-18
c3702 n10__i13__net7 vss 40.9884e-18
c3703 n5__r0_buff vss 63.9214e-18
c3704 n5__r1_buff vss 69.925e-18
c3705 n5__r2_buff vss 67.2136e-18
c3706 n8__i13__i19__net1 vss 63.5072e-18
c3707 n8__i13__i18__net1 vss 63.3692e-18
c3708 n7__i2__net1 vss 113.495e-18
c3709 n7__i1__net1 vss 117.079e-18
c3710 n7__i0__net1 vss 111.833e-18
c3711 n677__i18__net5 vss 596.013e-18
c3712 n5__net4 vss 90.4037e-18
c3713 n5__net3 vss 94.4327e-18
c3714 n6__i2__net79 vss 52.8263e-18
c3715 n6__i1__net79 vss 55.0232e-18
c3716 n6__i0__net79 vss 52.913e-18
c3717 n658__i18__net5 vss 603.391e-18
c3718 n6__i9__i1__net1 vss 37.6921e-18
c3719 n13__i13__net12 vss 60.2329e-18
c3720 n18__i13__net2 vss 57.1734e-18
c3721 n3__i9__i1__net1 vss 54.857e-18
c3722 n645__i18__net5 vss 601.062e-18
c3723 n27__shift vss 65.1545e-18
c3724 n13__reset_buff vss 64.3282e-18
c3725 n9__i13__net12 vss 105.368e-18
c3726 n11__i13__net2 vss 103.561e-18
c3727 n20__i13__a3 vss 89.1905e-18
c3728 n20__i13__a1 vss 88.8774e-18
c3729 n10__reset_buff vss 72.7892e-18
c3730 n638__i18__net5 vss 602.195e-18
c3731 n3__i13__i17__i4__net2 vss 23.4467e-18
c3732 n5__i13__i16__i4__net2 vss 2.77664e-18
c3733 n9__i9__net1 vss 50.6642e-18
c3734 n26__ck_buff vss 48.5609e-18
c3735 n80__vdd vss 74.3855e-18
c3736 n79__vdd vss 74.4032e-18
c3737 n227__vdd vss 88.9626e-18
c3738 n576__vddio vss 462.912e-18
c3739 n228__vdd vss 104.649e-18
c3740 n13__net14 vss 47.1117e-18
c3741 n8__i9__net2 vss 57.1382e-18
c3742 n15__ck_buff vss 69.9405e-18
c3743 n378__vdd vss 45.0147e-18
c3744 n12__i13__net11 vss 72.9422e-18
c3745 n14__i13__net1 vss 72.9583e-18
c3746 n624__i18__net5 vss 832.102e-18
c3747 n229__vdd vss 64.1955e-18
c3748 n24__ck_buff vss 57.6945e-18
c3749 n11__net14 vss 28.7528e-18
c3750 n6__i9__net2 vss 51.0757e-18
c3751 n13__ck_buff vss 75.4031e-18
c3752 n10__i13__net11 vss 41.0056e-18
c3753 n12__i13__net1 vss 40.9055e-18
c3754 n619__i18__net5 vss 462.842e-18
c3755 n230__vdd vss 79.4882e-18
c3756 n82__vdd vss 70.6535e-18
c3757 n81__vdd vss 70.6535e-18
c3758 n580__vddio vss 462.764e-18
c3759 n231__vdd vss 57.2608e-18
c3760 n10__i13__i17__net1 vss 77.3118e-18
c3761 n10__i13__i16__net1 vss 77.309e-18
c3762 n379__vdd vss 36.5415e-18
c3763 n13__net13 vss 49.1078e-18
c3764 n10__i9__i4__net4 vss 45.547e-18
c3765 n84__vdd vss 57.3481e-18
c3766 n83__vdd vss 57.3544e-18
c3767 n13__net10 vss 44.7973e-18
c3768 n611__i18__net5 vss 832.122e-18
c3769 n232__vdd vss 52.6491e-18
c3770 n233__vdd vss 84.6555e-18
c3771 n8__i13__i17__net1 vss 60.0128e-18
c3772 n8__i13__i16__net1 vss 62.1928e-18
c3773 n14__net13 vss 29.4343e-18
c3774 n8__i9__i4__net4 vss 60.3848e-18
c3775 n11__net10 vss 29.189e-18
c3776 n606__i18__net5 vss 602.583e-18
c3777 n584__vddio vss 462.602e-18
c3778 n380__vdd vss 53.4705e-18
c3779 n234__vdd vss 26.4334e-18
c3780 n16__net12 vss 56.9722e-18
c3781 n603__i18__net5 vss 828.563e-18
c3782 n13__net12 vss 35.8766e-18
c3783 n599__i18__net5 vss 530.211e-18
c3784 n381__vdd vss 62.899e-18
c3785 n235__vdd vss 51.2849e-18
c3786 n17__net12 vss 45.5535e-18
c3787 n614__vddio vss 416.593e-18
c3788 n14__i13__a3 vss 34.2927e-18
c3789 n13__i13__a1 vss 34.1761e-18
c3790 n9__i9__i4__net5 vss 38.132e-18
c3791 n21__x_out_3 vss 82.5055e-18
c3792 n22__x_out_1 vss 82.3954e-18
c3793 n382__vdd vss 75.5921e-18
c3794 n585__i18__net5 vss 855.309e-18
c3795 n13__i9__i4__net5 vss 84.7055e-18
c3796 n12__reset_b vss 69.1894e-18
c3797 n6__i9__i4__net2 vss 86.2954e-18
c3798 n10__i13__a3 vss 647.481e-21
c3799 n10__i13__a1 vss 647.481e-21
c3800 n18__net12 vss 31.7187e-18
c3801 n13__i13__a3 vss 51.6035e-18
c3802 n16__i13__a1 vss 50.2003e-18
c3803 n8__i9__i4__net5 vss 39.272e-18
c3804 n10__i13__i15__net2 vss 43.3004e-21
c3805 n8__i13__i13__net2 vss 43.4226e-21
c3806 n580__i18__net5 vss 469.392e-18
c3807 n12__i9__i4__net5 vss 62.4968e-18
c3808 n10__reset_b vss 69.9803e-18
c3809 n10__i9__i4__net2 vss 36.6193e-18
c3810 n9__i13__a3 vss 106.211e-18
c3811 n9__i13__a1 vss 113.345e-18
c3812 n383__vdd vss 104.144e-18
c3813 n617__vddio vss 416.591e-18
c3814 n15__y_out_3 vss 82.4295e-21
c3815 n236__vdd vss 92.816e-18
c3816 n9__reset_b vss 47.7991e-18
c3817 n237__vdd vss 47.3568e-18
c3818 n11__i9__i4__net2 vss 48.0118e-18
c3819 n5__i13__i15__net2 vss 110.858e-18
c3820 n3__i13__i13__net2 vss 110.394e-18
c3821 n572__i18__net5 vss 854.769e-18
c3822 n13__net9 vss 42.4772e-18
c3823 n238__vdd vss 98.0608e-18
c3824 n86__vdd vss 66.983e-18
c3825 n85__vdd vss 66.1696e-18
c3826 n13__y_out_3 vss 89.4003e-18
c3827 n12__y_out_1 vss 91.0374e-18
c3828 n7__reset_b vss 62.7413e-18
c3829 n9__i9__i4__net2 vss 60.4161e-18
c3830 n3__i13__i15__net2 vss 21.211e-18
c3831 n5__i13__i13__net2 vss 31.0602e-21
c3832 n567__i18__net5 vss 613.453e-18
c3833 n11__net9 vss 25.1981e-18
c3834 n590__vddio vss 462.879e-18
c3835 n564__i18__net5 vss 836.415e-18
c3836 n239__vdd vss 51.5424e-18
c3837 n16__net11 vss 58.1716e-18
c3838 n594__vddio vss 462.753e-18
c3839 n15__i9__i4__net1 vss 64.5845e-18
c3840 n560__i18__net5 vss 607.982e-18
c3841 n13__net11 vss 31.1509e-18
c3842 n240__vdd vss 64.0037e-18
c3843 n16__i13__a2 vss 39.0129e-18
c3844 n15__i13__a0 vss 36.0741e-18
c3845 n241__vdd vss 94.5634e-18
c3846 n17__net11 vss 46.2702e-18
c3847 n22__x_out_2 vss 81.4074e-18
c3848 n18__y_out_0 vss 81.4497e-18
c3849 n546__i18__net5 vss 832.166e-18
c3850 n9__i9__i4__net1 vss 41.526e-18
c3851 n10__i13__a2 vss 36.7693e-21
c3852 n10__i13__a0 vss 36.7693e-21
c3853 n242__vdd vss 78.687e-18
c3854 n598__vddio vss 462.611e-18
c3855 n11__ck_b vss 69.0427e-18
c3856 n13__i9__i4__net1 vss 90.8401e-18
c3857 n6__ck4 vss 51.386e-18
c3858 n15__i13__a2 vss 52.1634e-18
c3859 n18__i13__a0 vss 50.8786e-18
c3860 n18__net11 vss 28.3279e-18
c3861 n541__i18__net5 vss 602.539e-18
c3862 n8__i9__i4__net1 vss 36.0252e-18
c3863 n9__i13__a2 vss 105.029e-18
c3864 n9__i13__a0 vss 105.787e-18
c3865 n12__y_out_2 vss 86.7692e-18
c3866 n14__x_out_0 vss 90.2997e-18
c3867 n9__ck_b vss 75.7268e-18
c3868 n12__i9__i4__net1 vss 57.2936e-18
c3869 n8__ck4 vss 51.0112e-18
c3870 n528__i18__net5 vss 594.484e-18
c3871 n3__i13__i14__net2 vss 22.2357e-18
c3872 n243__vdd vss 108.564e-18
c3873 n533__i18__net5 vss 825.254e-18
c3874 n5__i13__i14__net2 vss 113.003e-18
c3875 n3__i13__i12__net2 vss 113.455e-18
c3876 n5__ck_b vss 65.7331e-18
c3877 n7__ck_b vss 55.8842e-18
c3878 n88__vdd vss 74.702e-18
c3879 n87__vdd vss 74.8815e-18
c3880 n602__vddio vss 462.655e-18
c3881 n245__vdd vss 74.1983e-18
c3882 n244__vdd vss 72.1406e-18
c3883 n9__y_out_3 vss 81.6167e-18
c3884 n7__y_out_2 vss 79.9415e-18
c3885 n9__y_out_1 vss 91.5859e-18
c3886 n9__y_out_0 vss 89.7644e-18
c3887 n520__i18__net5 vss 831.168e-18
c3888 n94__i14__net9 vss 68.5092e-18
c3889 n103__i14__net10 vss 122.073e-18
c3890 n385__vdd vss 90.7205e-18
c3891 n384__vdd vss 90.4268e-18
c3892 n90__vdd vss 90.8937e-18
c3893 n89__vdd vss 91.5324e-18
c3894 n606__vddio vss 464.299e-18
c3895 n247__vdd vss 108.472e-18
c3896 n246__vdd vss 105.299e-18
c3897 n9__i14__x_out_b_1 vss 57.7119e-18
c3898 n10__i14__y_out_b_2 vss 57.7635e-18
c3899 n9__i14__y_out_b_1 vss 57.7962e-18
c3900 n10__i14__x_out_b_0 vss 57.8044e-18
c3901 n91__i14__net9 vss 68.2144e-18
c3902 n100__i14__net10 vss 122.844e-18
c3903 n387__vdd vss 64.9258e-18
c3904 n386__vdd vss 64.7769e-18
c3905 n92__vdd vss 64.7881e-18
c3906 n91__vdd vss 64.8394e-18
c3907 n510__i18__net5 vss 844.488e-18
c3908 n249__vdd vss 108.46e-18
c3909 n248__vdd vss 103.482e-18
c3910 n389__vdd vss 58.554e-18
c3911 n388__vdd vss 58.5707e-18
c3912 n94__vdd vss 58.6124e-18
c3913 n93__vdd vss 58.6522e-18
c3914 n88__i14__net9 vss 67.7631e-18
c3915 n97__i14__net10 vss 117.871e-18
c3916 n610__vddio vss 258.361e-18
c3917 n11__i14__i11__net4 vss 46.4831e-18
c3918 n11__i14__i14__net4 vss 46.3698e-18
c3919 n11__i14__i15__net4 vss 46.468e-18
c3920 n11__i14__i12__net4 vss 46.3852e-18
c3921 n251__vdd vss 90.4804e-18
c3922 n250__vdd vss 50.8989e-18
c3923 n391__vdd vss 92.3563e-18
c3924 n390__vdd vss 92.4655e-18
c3925 n96__vdd vss 92.3433e-18
c3926 n95__vdd vss 92.462e-18
c3927 n252__vdd vss 52.2972e-18
c3928 n2__ck4 vss 55.2743e-18
c3929 n15__i14__i11__net5 vss 852.7e-21
c3930 n15__i14__i14__net5 vss 847.984e-21
c3931 n15__i14__i15__net5 vss 847.984e-21
c3932 n15__i14__i12__net5 vss 900.802e-21
c3933 n70__i14__net3 vss 116.578e-18
c3934 n253__vdd vss 110.611e-18
c3935 n393__vdd vss 27.032e-18
c3936 n392__vdd vss 26.8405e-18
c3937 n98__vdd vss 26.8455e-18
c3938 n97__vdd vss 26.5383e-18
c3939 n254__vdd vss 103.212e-18
c3940 n60__i14__net3 vss 127.345e-18
c3941 n395__vdd vss 52.3316e-18
c3942 n394__vdd vss 52.7696e-18
c3943 n100__vdd vss 52.6878e-18
c3944 n99__vdd vss 52.5374e-18
c3945 n255__vdd vss 58.1076e-18
c3946 n256__vdd vss 98.9446e-18
c3947 n9__i14__i11__net5 vss 40.7284e-18
c3948 n9__i14__i14__net5 vss 38.4224e-18
c3949 n9__i14__i15__net5 vss 40.7348e-18
c3950 n9__i14__i12__net5 vss 38.4224e-18
c3951 n57__i14__net3 vss 126.419e-18
c3952 n699__vddio vss 257.96e-18
c3953 n12__i14__i11__net5 vss 85.1966e-18
c3954 n13__i14__i14__net5 vss 85.2206e-18
c3955 n12__i14__i15__net5 vss 85.0628e-18
c3956 n13__i14__i12__net5 vss 85.2206e-18
c3957 n257__vdd vss 81.4251e-18
c3958 n258__vdd vss 61.9793e-18
c3959 n11__i14__i11__net2 vss 83.1632e-18
c3960 n6__i14__i14__net2 vss 82.9699e-18
c3961 n11__i14__i15__net2 vss 83.1632e-18
c3962 n6__i14__i12__net2 vss 82.9699e-18
c3963 n648__r_out vss 895.064e-18
c3964 n57__i14__net4 vss 69.7043e-18
c3965 n397__vdd vss 93.5454e-18
c3966 n396__vdd vss 93.5963e-18
c3967 n102__vdd vss 93.5454e-18
c3968 n101__vdd vss 93.6768e-18
c3969 n18__i14__i17__net10 vss 68.2007e-18
c3970 n259__vdd vss 108.544e-18
c3971 n768__vddio vss 456.642e-18
c3972 n9__i14__i11__net2 vss 48.9651e-18
c3973 n11__i14__i14__net2 vss 48.8521e-18
c3974 n9__i14__i15__net2 vss 48.9651e-18
c3975 n11__i14__i12__net2 vss 48.8536e-18
c3976 n260__vdd vss 141.44e-18
c3977 n54__i14__net4 vss 69.188e-18
c3978 n399__vdd vss 97.3518e-18
c3979 n398__vdd vss 97.3291e-18
c3980 n104__vdd vss 97.3518e-18
c3981 n103__vdd vss 97.2979e-18
c3982 n264__vdd vss 110.388e-18
c3983 n263__vdd vss 141.409e-18
c3984 n635__r_out vss 958.265e-18
c3985 n51__i14__net4 vss 68.6191e-18
c3986 n18__i14__i17__net9 vss 115.24e-18
c3987 n772__vddio vss 455.276e-18
c3988 n265__vdd vss 84.2266e-18
c3989 n11__i14__i17__net10 vss 88.0222e-18
c3990 n266__vdd vss 115.935e-18
c3991 n25__i14__net7 vss 120.859e-18
c3992 n622__r_out vss 875.892e-18
c3993 n267__vdd vss 80.3158e-18
c3994 n268__vdd vss 118.963e-18
c3995 n401__vdd vss 93.826e-18
c3996 n400__vdd vss 93.8763e-18
c3997 n106__vdd vss 93.8763e-18
c3998 n105__vdd vss 93.8638e-18
c3999 n776__vddio vss 454.615e-18
c4000 n8__i14__i17__net9 vss 82.468e-18
c4001 n26__i14__net11 vss 52.8741e-18
c4002 n271__vdd vss 85.4434e-18
c4003 n9__i14__i11__net1 vss 40.8868e-18
c4004 n9__i14__i14__net1 vss 38.4504e-18
c4005 n9__i14__i15__net1 vss 40.8868e-18
c4006 n9__i14__i12__net1 vss 38.4504e-18
c4007 n609__r_out vss 880.758e-18
c4008 n12__i14__i11__net1 vss 88.6006e-18
c4009 n13__i14__i14__net1 vss 88.6331e-18
c4010 n12__i14__i15__net1 vss 88.6006e-18
c4011 n13__i14__i12__net1 vss 88.6331e-18
c4012 n19__i14__i17__net7 vss 86.9013e-18
c4013 n10__i14__i17__net11 vss 97.5495e-18
c4014 n780__vddio vss 454.523e-18
c4015 n3__y3 vss 56.6147e-18
c4016 n1__y2 vss 56.4406e-18
c4017 n3__y1 vss 56.6469e-18
c4018 n1__y0 vss 56.4406e-18
c4019 n273__vdd vss 87.8418e-18
c4020 n272__vdd vss 90.88e-18
c4021 n28__i14__i17__net1 vss 55.9625e-18
c4022 n22__i14__i17__net8 vss 57.8156e-18
c4023 n596__r_out vss 876.185e-18
c4024 n3__x_out_3 vss 97.5749e-18
c4025 n3__x_out_1 vss 97.5749e-18
c4026 n275__vdd vss 65.098e-18
c4027 n274__vdd vss 69.4993e-18
c4028 n403__vdd vss 94.9481e-18
c4029 n402__vdd vss 94.9481e-18
c4030 n108__vdd vss 94.9481e-18
c4031 n107__vdd vss 94.8852e-18
c4032 n784__vddio vss 454.383e-18
c4033 n277__vdd vss 58.5985e-18
c4034 n276__vdd vss 60.8526e-18
c4035 n9__i14__y_out_b_3 vss 58.1119e-18
c4036 n10__i14__y_out_b_0 vss 58.1312e-18
c4037 n9__i14__x_out_b_2 vss 58.1312e-18
c4038 n10__i14__x_out_b_3 vss 58.1312e-18
c4039 n10__i14__i17__i2__net4 vss 45.6508e-18
c4040 n10__i14__i17__i3__net4 vss 44.6588e-18
c4041 n405__vdd vss 64.7569e-18
c4042 n404__vdd vss 64.6924e-18
c4043 n110__vdd vss 64.6924e-18
c4044 n109__vdd vss 64.6924e-18
c4045 n583__r_out vss 881.273e-18
c4046 n279__vdd vss 92.625e-18
c4047 n278__vdd vss 94.3993e-18
c4048 n407__vdd vss 58.647e-18
c4049 n406__vdd vss 58.6636e-18
c4050 n112__vdd vss 58.6636e-18
c4051 n111__vdd vss 58.7626e-18
c4052 n788__vddio vss 454.573e-18
c4053 n10__i14__i13__net4 vss 46.8414e-18
c4054 n10__i14__i16__net4 vss 46.6871e-18
c4055 n10__i14__i10__net4 vss 46.8052e-18
c4056 n10__i14__i9__net4 vss 46.6755e-18
c4057 n15__i14__i17__i2__net5 vss 16.8525e-21
c4058 n281__vdd vss 26.5821e-18
c4059 n280__vdd vss 26.7512e-18
c4060 n409__vdd vss 92.4637e-18
c4061 n408__vdd vss 92.2466e-18
c4062 n114__vdd vss 92.476e-18
c4063 n113__vdd vss 92.2466e-18
c4064 n570__r_out vss 877.158e-18
c4065 n283__vdd vss 51.4446e-18
c4066 n282__vdd vss 50.9502e-18
c4067 n792__vddio vss 454.016e-18
c4068 n411__vdd vss 25.9672e-18
c4069 n410__vdd vss 25.5735e-18
c4070 n116__vdd vss 25.8451e-18
c4071 n115__vdd vss 25.1809e-18
c4072 n9__i14__i17__i2__net5 vss 40.4858e-18
c4073 n9__i14__i17__i3__net5 vss 38.2536e-18
c4074 n413__vdd vss 50.3283e-18
c4075 n412__vdd vss 51.0274e-18
c4076 n120__vdd vss 51.0274e-18
c4077 n117__vdd vss 50.5488e-18
c4078 n557__r_out vss 878.698e-18
c4079 n12__i14__i17__i2__net5 vss 85.5842e-18
c4080 n13__i14__i17__i3__net5 vss 85.8352e-18
c4081 n11__i14__i17__i2__net2 vss 82.4252e-18
c4082 n6__i14__i17__i3__net2 vss 81.8663e-18
c4083 n9__i14__i13__net5 vss 42.1669e-18
c4084 n9__i14__i16__net5 vss 39.7124e-18
c4085 n9__i14__i10__net5 vss 42.1645e-18
c4086 n9__i14__i9__net5 vss 39.7124e-18
c4087 n796__vddio vss 453.649e-18
c4088 n285__vdd vss 92.5109e-18
c4089 n284__vdd vss 93.9092e-18
c4090 n12__i14__i13__net5 vss 84.5514e-18
c4091 n13__i14__i16__net5 vss 84.6372e-18
c4092 n12__i14__i10__net5 vss 84.7369e-18
c4093 n13__i14__i9__net5 vss 84.7694e-18
c4094 n544__r_out vss 874.232e-18
c4095 n9__i14__i17__i2__net2 vss 47.5296e-18
c4096 n11__i14__i17__i3__net2 vss 48.2315e-18
c4097 n11__i14__i13__net2 vss 82.2903e-18
c4098 n6__i14__i16__net2 vss 82.0671e-18
c4099 n11__i14__i10__net2 vss 82.2903e-18
c4100 n6__i14__i9__net2 vss 82.0671e-18
c4101 n287__vdd vss 96.6575e-18
c4102 n286__vdd vss 97.6975e-18
c4103 n415__vdd vss 92.6636e-18
c4104 n414__vdd vss 92.8729e-18
c4105 n123__vdd vss 92.6728e-18
c4106 n119__vdd vss 92.8729e-18
c4107 n800__vddio vss 455.013e-18
c4108 n9__i14__i13__net2 vss 48.7405e-18
c4109 n11__i14__i16__net2 vss 48.6275e-18
c4110 n9__i14__i10__net2 vss 48.7405e-18
c4111 n11__i14__i9__net2 vss 48.6275e-18
c4112 n531__r_out vss 879.021e-18
c4113 n417__vdd vss 97.6267e-18
c4114 n416__vdd vss 97.6267e-18
c4115 n127__vdd vss 97.6267e-18
c4116 n122__vdd vss 97.6267e-18
c4117 n804__vddio vss 454.546e-18
c4118 n289__vdd vss 94.5989e-18
c4119 n288__vdd vss 93.8933e-18
c4120 n521__r_out vss 877.584e-18
c4121 n9__i14__i17__i2__net1 vss 40.8504e-18
c4122 n9__i14__i17__i3__net1 vss 38.187e-18
c4123 n808__vddio vss 453.552e-18
c4124 n418__vdd vss 95.1363e-18
c4125 n348__vdd vss 95.3333e-18
c4126 n129__vdd vss 95.3333e-18
c4127 n126__vdd vss 95.1814e-18
c4128 n12__i14__i17__i2__net1 vss 88.779e-18
c4129 n13__i14__i17__i3__net1 vss 88.0621e-18
c4130 n510__r_out vss 871.492e-18
c4131 n7__i14__i17__net1 vss 58.529e-18
c4132 n9__i14__i13__net1 vss 41.8275e-18
c4133 n9__i14__i16__net1 vss 39.4826e-18
c4134 n9__i14__i10__net1 vss 41.9078e-18
c4135 n9__i14__i9__net1 vss 39.4703e-18
c4136 n812__vddio vss 453.973e-18
c4137 n7__i14__i17__net3 vss 81.231e-18
c4138 n5__i14__i17__net6 vss 93.6712e-18
c4139 n12__i14__i13__net1 vss 88.9635e-18
c4140 n13__i14__i16__net1 vss 89.0013e-18
c4141 n12__i14__i10__net1 vss 88.8198e-18
c4142 n13__i14__i9__net1 vss 88.8519e-18
c4143 n290__vdd vss 45.7251e-18
c4144 n210__vdd vss 37.8168e-18
c4145 n3__x3 vss 54.6354e-18
c4146 n1__x2 vss 54.4405e-18
c4147 n3__x1 vss 54.6354e-18
c4148 n1__x0 vss 54.4405e-18
c4149 n7__y_out_3 vss 45.2373e-18
c4150 n9__y_out_2 vss 42.9906e-18
c4151 n7__y_out_1 vss 50.7784e-18
c4152 n11__y_out_0 vss 52.5598e-18
c4153 n515__i18__net5 vss 648.665e-18
c4154 n92__i14__net9 vss 77.8166e-18
c4155 n105__i14__net10 vss 79.5069e-18
c4156 n10__i14__x_out_b_1 vss 58.6221e-18
c4157 n8__i14__y_out_b_2 vss 50.8309e-18
c4158 n10__i14__y_out_b_1 vss 51.1218e-18
c4159 n8__i14__x_out_b_0 vss 51.3301e-18
c4160 n89__i14__net9 vss 80.8819e-18
c4161 n102__i14__net10 vss 88.6448e-18
c4162 n506__i18__net5 vss 611.8e-18
c4163 n86__i14__net9 vss 78.3989e-18
c4164 n99__i14__net10 vss 81.768e-18
c4165 n9__i14__i11__net4 vss 67.291e-18
c4166 n9__i14__i14__net4 vss 63.3142e-18
c4167 n9__i14__i15__net4 vss 63.2873e-18
c4168 n9__i14__i12__net4 vss 62.2132e-18
c4169 n71__i14__net3 vss 79.2908e-18
c4170 n2__i14__clk_div4_out_b vss 6.48822e-21
c4171 n62__i14__net3 vss 91.0294e-18
c4172 n8__i14__i11__net5 vss 37.9702e-18
c4173 n8__i14__i14__net5 vss 36.9733e-18
c4174 n8__i14__i15__net5 vss 34.6431e-18
c4175 n8__i14__i12__net5 vss 38.2888e-18
c4176 n59__i14__net3 vss 83.6691e-18
c4177 n13__i14__i11__net5 vss 58.5319e-18
c4178 n12__i14__i14__net5 vss 55.4318e-18
c4179 n13__i14__i15__net5 vss 55.5105e-18
c4180 n12__i14__i12__net5 vss 59.7545e-18
c4181 n6__i14__i11__net2 vss 37.1576e-18
c4182 n10__i14__i14__net2 vss 35.1566e-18
c4183 n6__i14__i15__net2 vss 35.068e-18
c4184 n10__i14__i12__net2 vss 37.918e-18
c4185 n643__r_out vss 516.23e-18
c4186 n55__i14__net4 vss 80.0717e-18
c4187 n20__i14__i17__net10 vss 48.1563e-18
c4188 n12__i14__i11__net2 vss 59.0767e-18
c4189 n9__i14__i14__net2 vss 58.861e-18
c4190 n12__i14__i15__net2 vss 58.8891e-18
c4191 n9__i14__i12__net2 vss 60.5977e-18
c4192 n262__vdd vss 94.9089e-18
c4193 n52__i14__net4 vss 82.7495e-18
c4194 n630__r_out vss 643.886e-18
c4195 n49__i14__net4 vss 80.7251e-18
c4196 n20__i14__i17__net9 vss 52.2817e-18
c4197 n15__i14__i11__net1 vss 67.9386e-18
c4198 n15__i14__i14__net1 vss 65.2865e-18
c4199 n15__i14__i15__net1 vss 65.2674e-18
c4200 n15__i14__i12__net1 vss 64.0433e-18
c4201 n13__i14__i17__net10 vss 74.4763e-18
c4202 n617__r_out vss 505.449e-18
c4203 n270__vdd vss 107.869e-18
c4204 n10__i14__i17__net9 vss 29.8085e-18
c4205 n25__i14__net11 vss 114.493e-18
c4206 n8__i14__i11__net1 vss 36.1897e-18
c4207 n8__i14__i14__net1 vss 35.9321e-18
c4208 n8__i14__i15__net1 vss 33.7432e-18
c4209 n8__i14__i12__net1 vss 36.1695e-18
c4210 n604__r_out vss 509.976e-18
c4211 n13__i14__i11__net1 vss 60.4935e-18
c4212 n12__i14__i14__net1 vss 56.4676e-18
c4213 n13__i14__i15__net1 vss 56.5177e-18
c4214 n12__i14__i12__net1 vss 57.1923e-18
c4215 n17__i14__i17__net7 vss 51.893e-18
c4216 n12__i14__i17__net11 vss 50.3194e-18
c4217 n1__y3 vss 58.1063e-18
c4218 n3__y2 vss 58.0174e-18
c4219 n1__y1 vss 57.8861e-18
c4220 n3__y0 vss 58.106e-18
c4221 n29__i14__i17__net1 vss 47.9435e-18
c4222 n20__i14__i17__net8 vss 48.7229e-18
c4223 n591__r_out vss 646.736e-18
c4224 n3__x_out_2 vss 56.2792e-18
c4225 n3__x_out_0 vss 56.8214e-18
c4226 n10__i14__y_out_b_3 vss 60.0689e-18
c4227 n8__i14__y_out_b_0 vss 53.2552e-18
c4228 n10__i14__x_out_b_2 vss 53.2552e-18
c4229 n8__i14__x_out_b_3 vss 56.0372e-18
c4230 n8__i14__i17__i2__net4 vss 64.7735e-18
c4231 n8__i14__i17__i3__net4 vss 64.9824e-18
c4232 n578__r_out vss 506.733e-18
c4233 n8__i14__i13__net4 vss 68.7973e-18
c4234 n8__i14__i16__net4 vss 62.9844e-18
c4235 n8__i14__i10__net4 vss 62.9844e-18
c4236 n8__i14__i9__net4 vss 64.8953e-18
c4237 n565__r_out vss 580.492e-18
c4238 n8__i14__i17__i2__net5 vss 34.2581e-18
c4239 n8__i14__i17__i3__net5 vss 37.3557e-18
c4240 n552__r_out vss 578.285e-18
c4241 n13__i14__i17__i2__net5 vss 54.7286e-18
c4242 n12__i14__i17__i3__net5 vss 55.5788e-18
c4243 n6__i14__i17__i2__net2 vss 33.6493e-18
c4244 n10__i14__i17__i3__net2 vss 34.6666e-18
c4245 n8__i14__i13__net5 vss 33.194e-18
c4246 n8__i14__i16__net5 vss 35.4501e-18
c4247 n8__i14__i10__net5 vss 33.1914e-18
c4248 n8__i14__i9__net5 vss 36.4331e-18
c4249 n13__i14__i13__net5 vss 56.8747e-18
c4250 n12__i14__i16__net5 vss 54.357e-18
c4251 n13__i14__i10__net5 vss 53.8936e-18
c4252 n12__i14__i9__net5 vss 56.0043e-18
c4253 n539__r_out vss 503.628e-18
c4254 n12__i14__i17__i2__net2 vss 59.1408e-18
c4255 n9__i14__i17__i3__net2 vss 61.6453e-18
c4256 n6__i14__i13__net2 vss 34.2744e-18
c4257 n10__i14__i16__net2 vss 33.5806e-18
c4258 n6__i14__i10__net2 vss 33.483e-18
c4259 n10__i14__i9__net2 vss 34.528e-18
c4260 n12__i14__i13__net2 vss 61.0109e-18
c4261 n9__i14__i16__net2 vss 60.2079e-18
c4262 n12__i14__i10__net2 vss 60.2323e-18
c4263 n9__i14__i9__net2 vss 63.0706e-18
c4264 n526__r_out vss 586.415e-18
c4265 n15__i14__i17__i2__net1 vss 63.4567e-18
c4266 n15__i14__i17__i3__net1 vss 64.6289e-18
c4267 n15__i14__i13__net1 vss 65.6221e-18
c4268 n15__i14__i16__net1 vss 65.0118e-18
c4269 n15__i14__i10__net1 vss 64.9926e-18
c4270 n15__i14__i9__net1 vss 65.8741e-18
c4271 n517__r_out vss 508.794e-18
c4272 n8__i14__i17__i2__net1 vss 33.0581e-18
c4273 n8__i14__i17__i3__net1 vss 37.2295e-18
c4274 n13__i14__i17__i2__net1 vss 55.6957e-18
c4275 n12__i14__i17__i3__net1 vss 57.9753e-18
c4276 n506__r_out vss 645.585e-18
c4277 n5__i14__i17__net1 vss 59.4687e-18
c4278 n3__i14__i17__net8 vss 65.2319e-18
c4279 n8__i14__i13__net1 vss 33.8638e-18
c4280 n8__i14__i16__net1 vss 35.6146e-18
c4281 n8__i14__i10__net1 vss 33.4512e-18
c4282 n8__i14__i9__net1 vss 37.3218e-18
c4283 n5__i14__i17__net3 vss 52.6118e-18
c4284 n7__i14__i17__net6 vss 39.0659e-18
c4285 n13__i14__i13__net1 vss 58.1051e-18
c4286 n12__i14__i16__net1 vss 58.1574e-18
c4287 n13__i14__i10__net1 vss 58.1712e-18
c4288 n12__i14__i9__net1 vss 58.6823e-18
c4289 n1__x3 vss 50.7257e-18
c4290 n3__x2 vss 50.3508e-18
c4291 n1__x1 vss 50.1882e-18
c4292 n3__x0 vss 52.4004e-18
c4293 n497__r_out vss 878.042e-18
c4294 n816__vddio vss 454.615e-18
c4295 n482__r_out vss 878.714e-18
c4296 n820__vddio vss 454.523e-18
c4297 n466__r_out vss 877.099e-18
c4298 n824__vddio vss 453.675e-18
c4299 n450__r_out vss 876.055e-18
c4300 n828__vddio vss 453.558e-18
c4301 n442__r_out vss 869.281e-18
c4302 n832__vddio vss 455.408e-18
c4303 n422__r_out vss 881.497e-18
c4304 n836__vddio vss 455.078e-18
c4305 n409__r_out vss 877.578e-18
c4306 n840__vddio vss 453.54e-18
c4307 n399__r_out vss 875.561e-18
c4308 n844__vddio vss 454.953e-18
c4309 n386__r_out vss 878.714e-18
c4310 n848__vddio vss 454.541e-18
c4311 n375__r_out vss 877.099e-18
c4312 n852__vddio vss 453.942e-18
c4313 n360__r_out vss 876.056e-18
c4314 n856__vddio vss 453.596e-18
c4315 n344__r_out vss 871.72e-18
c4316 n860__vddio vss 454.981e-18
c4317 n336__r_out vss 879.018e-18
c4318 n864__vddio vss 455.83e-18
c4319 n323__r_out vss 877.578e-18
c4320 n868__vddio vss 453.558e-18
c4321 n310__r_out vss 871.495e-18
c4322 n872__vddio vss 453.962e-18
c4323 n297__r_out vss 878.093e-18
c4324 n876__vddio vss 454.62e-18
c4325 n279__r_out vss 878.652e-18
c4326 n880__vddio vss 454.529e-18
c4327 n271__r_out vss 877.102e-18
c4328 n884__vddio vss 453.817e-18
c4329 n258__r_out vss 876.11e-18
c4330 n888__vddio vss 453.558e-18
c4331 n245__r_out vss 861.744e-18
c4332 n892__vddio vss 448.312e-18
c4333 n232__r_out vss 864.315e-18
c4334 n896__vddio vss 447.87e-18
c4335 n214__r_out vss 860.435e-18
c4336 n900__vddio vss 446.207e-18
c4337 n206__r_out vss 860.643e-18
c4338 n904__vddio vss 447.87e-18
c4339 n191__r_out vss 851.597e-18
c4340 n908__vddio vss 452.086e-18
c4341 n180__r_out vss 860.059e-18
c4342 n912__vddio vss 448.151e-18
c4343 n165__r_out vss 862.125e-18
c4344 n916__vddio vss 451.078e-18
c4345 n149__r_out vss 858.648e-18
c4346 n920__vddio vss 447.178e-18
c4347 n136__r_out vss 863.477e-18
c4348 n924__vddio vss 447.318e-18
c4349 n128__r_out vss 875.213e-18
c4350 n928__vddio vss 453.555e-18
c4351 n115__r_out vss 868.691e-18
c4352 n932__vddio vss 445.997e-18
c4353 n102__r_out vss 853.058e-18
c4354 n936__vddio vss 447.816e-18
c4355 n84__r_out vss 854.77e-18
c4356 n940__vddio vss 447.724e-18
c4357 n76__r_out vss 858.694e-18
c4358 n944__vddio vss 448.297e-18
c4359 n61__r_out vss 859.416e-18
c4360 n948__vddio vss 448.386e-18
c4361 n50__r_out vss 855.989e-18
c4362 n952__vddio vss 447.927e-18
c4363 n35__r_out vss 860.955e-18
c4364 n493__r_out vss 578.748e-18
c4365 n478__r_out vss 506.101e-18
c4366 n461__r_out vss 647.279e-18
c4367 n445__r_out vss 642.929e-18
c4368 n438__r_out vss 639.642e-18
c4369 n417__r_out vss 649.424e-18
c4370 n404__r_out vss 644.68e-18
c4371 n395__r_out vss 645.78e-18
c4372 n382__r_out vss 505.952e-18
c4373 n371__r_out vss 647.092e-18
c4374 n356__r_out vss 504.131e-18
c4375 n339__r_out vss 499.489e-18
c4376 n332__r_out vss 649.656e-18
c4377 n319__r_out vss 644.68e-18
c4378 n306__r_out vss 641.722e-18
c4379 n293__r_out vss 645.611e-18
c4380 n274__r_out vss 645.304e-18
c4381 n267__r_out vss 646.984e-18
c4382 n254__r_out vss 642.888e-18
c4383 n241__r_out vss 639.642e-18
c4384 n228__r_out vss 649.477e-18
c4385 n209__r_out vss 644.627e-18
c4386 n202__r_out vss 644.959e-18
c4387 n187__r_out vss 501.19e-18
c4388 n176__r_out vss 645.765e-18
c4389 n161__r_out vss 506.226e-18
c4390 n144__r_out vss 503.198e-18
c4391 n131__r_out vss 648.99e-18
c4392 n124__r_out vss 645.726e-18
c4393 n111__r_out vss 640.166e-18
c4394 n98__r_out vss 630.581e-18
c4395 n79__r_out vss 630.179e-18
c4396 n72__r_out vss 635.984e-18
c4397 n57__r_out vss 496.352e-18
c4398 n46__r_out vss 634.107e-18
c4399 n31__r_out vss 498.606e-18
c4400 n14__r_out vss 496.825e-18
c4401 n7__r_out vss 641.117e-18
c4402 n956__vddio vss 447.575e-18
c4403 n19__r_out vss 859.841e-18
c4404 n960__vddio vss 447.345e-18
c4405 n11__r_out vss 864.134e-18
c4406 n762__vddio vss 266.299e-18
c4407 n2__i14__i13__net1 vss 16.8064e-18
c4408 n3__i14__i13__net1 vss 8.85348e-18
c4409 n2__i14__i16__net1 vss 16.4865e-18
c4410 n3__i14__i16__net1 vss 8.84604e-18
c4411 n2__i14__i10__net1 vss 18.8428e-18
c4412 n3__i14__i10__net1 vss 10.5544e-18
c4413 n2__i14__i9__net1 vss 17.6041e-18
c4414 n3__i14__i9__net1 vss 8.5021e-18
c4415 n2__i14__i17__i2__net1 vss 16.3128e-18
c4416 n3__i14__i17__i2__net1 vss 8.00073e-18
c4417 n2__i14__i17__i3__net1 vss 15.7708e-18
c4418 n3__i14__i17__i3__net1 vss 8.30759e-18
c4419 n2__i14__i13__net5 vss 18.611e-18
c4420 n3__i14__i13__net5 vss 12.3122e-18
c4421 n2__i14__i16__net5 vss 19.0843e-18
c4422 n3__i14__i16__net5 vss 10.2793e-18
c4423 n2__i14__i10__net5 vss 19.7326e-18
c4424 n3__i14__i10__net5 vss 11.9836e-18
c4425 n2__i14__i9__net5 vss 18.1396e-18
c4426 n3__i14__i9__net5 vss 9.38222e-18
c4427 n2__i14__i17__i2__net5 vss 17.0944e-18
c4428 n3__i14__i17__i2__net5 vss 9.02404e-18
c4429 n2__i14__i17__i3__net5 vss 17.588e-18
c4430 n3__i14__i17__i3__net5 vss 9.15435e-18
c4431 n9__ck vss 29.2943e-18
c4432 n10__ck vss 36.0674e-18
c4433 n9__reset vss 18.1219e-18
c4434 n10__reset vss 35.7765e-18
c4435 n17__i14__net10 vss 34.2747e-18
c4436 n19__i14__net10 vss 54.984e-18
c4437 n20__i14__net10 vss 55.131e-18
c4438 n21__i14__net10 vss 34.0171e-18
c4439 n23__i14__net10 vss 34.2747e-18
c4440 n25__i14__net10 vss 54.9905e-18
c4441 n26__i14__net10 vss 55.131e-18
c4442 n27__i14__net10 vss 34.0171e-18
c4443 n2__i14__y_out_b_3 vss 11.3986e-18
c4444 n2__i14__y_out_b_0 vss 10.1258e-18
c4445 n2__i14__x_out_b_2 vss 9.60454e-18
c4446 n2__i14__x_out_b_3 vss 10.1258e-18
c4447 n12__ck vss 34.8367e-18
c4448 n14__ck vss 54.9729e-18
c4449 n5__i14__i17__net7 vss 55.4793e-18
c4450 n6__i14__i17__net7 vss 34.5791e-18
c4451 n15__i14__i17__net1 vss 10.4223e-18
c4452 n7__i14__i17__net8 vss 9.11932e-18
c4453 n2__i14__i17__net10 vss 10.6977e-18
c4454 n21__i14__net3 vss 46.6779e-18
c4455 n22__i14__net3 vss 47.4625e-18
c4456 n23__i14__net3 vss 45.2798e-18
c4457 n24__i14__net3 vss 46.3923e-18
c4458 n25__i14__net3 vss 46.6779e-18
c4459 n26__i14__net3 vss 44.9889e-18
c4460 n27__i14__net3 vss 44.8731e-18
c4461 n2__i14__i17__net9 vss 11.3946e-18
c4462 n16__reset vss 46.5216e-18
c4463 n18__reset vss 44.0189e-18
c4464 n20__reset vss 44.8696e-18
c4465 n21__reset vss 48.1344e-18
c4466 n7__i14__i13__net2 vss 91.9212e-18
c4467 n8__i14__i13__net2 vss 59.1425e-18
c4468 n7__i14__i16__net2 vss 91.3767e-18
c4469 n8__i14__i16__net2 vss 58.5975e-18
c4470 n7__i14__i10__net2 vss 90.8619e-18
c4471 n8__i14__i10__net2 vss 58.9312e-18
c4472 n7__i14__i9__net2 vss 91.1816e-18
c4473 n8__i14__i9__net2 vss 58.5388e-18
c4474 n2__i14__i11__net1 vss 17.2096e-18
c4475 n3__i14__i11__net1 vss 9.4067e-18
c4476 n2__i14__i14__net1 vss 16.9032e-18
c4477 n3__i14__i14__net1 vss 8.8989e-18
c4478 n2__i14__i15__net1 vss 17.2204e-18
c4479 n3__i14__i15__net1 vss 9.2441e-18
c4480 n2__i14__i12__net1 vss 15.5325e-18
c4481 n3__i14__i12__net1 vss 7.96158e-18
c4482 n7__i14__i17__i2__net2 vss 91.0893e-18
c4483 n8__i14__i17__i2__net2 vss 63.1105e-18
c4484 n7__i14__i17__i3__net2 vss 91.1875e-18
c4485 n8__i14__i17__i3__net2 vss 58.2481e-18
c4486 n27__reset vss 15.9201e-18
c4487 n28__reset vss 8.49841e-18
c4488 n30__reset vss 6.81903e-18
c4489 n31__reset vss 6.86627e-18
c4490 n33__reset vss 6.93013e-18
c4491 n34__reset vss 14.5181e-18
c4492 n2__i14__net7 vss 9.92452e-18
c4493 n2__i14__net11 vss 11.0013e-18
c4494 n30__i14__net4 vss 17.9823e-18
c4495 n31__i14__net4 vss 7.30446e-18
c4496 n33__i14__net4 vss 9.08929e-18
c4497 n34__i14__net4 vss 6.46747e-18
c4498 n36__i14__net4 vss 7.07438e-18
c4499 n37__i14__net4 vss 15.5257e-18
c4500 n2__i14__i11__net5 vss 20.4469e-18
c4501 n3__i14__i11__net5 vss 11.4054e-18
c4502 n2__i14__i14__net5 vss 19.3232e-18
c4503 n3__i14__i14__net5 vss 9.66976e-18
c4504 n2__i14__i15__net5 vss 18.8947e-18
c4505 n3__i14__i15__net5 vss 11.6769e-18
c4506 n2__i14__i12__net5 vss 18.9631e-18
c4507 n3__i14__i12__net5 vss 8.67291e-18
c4508 n7__i14__y_out_b_3 vss 45.4936e-18
c4509 n7__i14__y_out_b_0 vss 42.618e-18
c4510 n7__i14__x_out_b_2 vss 45.6427e-18
c4511 n7__i14__x_out_b_3 vss 42.618e-18
c4512 n26__i14__i17__net1 vss 41.0596e-18
c4513 n19__i14__i17__net8 vss 41.1952e-18
c4514 n65__i14__net10 vss 34.2747e-18
c4515 n67__i14__net10 vss 57.1751e-18
c4516 n68__i14__net10 vss 55.3833e-18
c4517 n69__i14__net10 vss 34.0171e-18
c4518 n71__i14__net10 vss 34.2747e-18
c4519 n73__i14__net10 vss 55.1364e-18
c4520 n74__i14__net10 vss 55.4431e-18
c4521 n75__i14__net10 vss 34.0171e-18
c4522 n31__i14__i17__net1 vss 32.1439e-18
c4523 n6__i14__net7 vss 14.0165e-18
c4524 n7__i14__net7 vss 6.88826e-18
c4525 n9__i14__net7 vss 6.76696e-18
c4526 n10__i14__net7 vss 6.8344e-18
c4527 n12__i14__net7 vss 7.0056e-18
c4528 n13__i14__net7 vss 15.3438e-18
c4529 n6__i14__net11 vss 13.8092e-18
c4530 n7__i14__net11 vss 6.81522e-18
c4531 n9__i14__net11 vss 7.22837e-18
c4532 n10__i14__net11 vss 6.66326e-18
c4533 n12__i14__net11 vss 8.26408e-18
c4534 n13__i14__net11 vss 17.3916e-18
c4535 n2__i14__x_out_b_1 vss 11.1097e-18
c4536 n2__i14__y_out_b_2 vss 9.3517e-18
c4537 n2__i14__y_out_b_1 vss 9.98756e-18
c4538 n2__i14__x_out_b_0 vss 9.93171e-18
c4539 n7__x_out_2 vss 8.86603e-18
c4540 n2__y_out_0 vss 8.31369e-18
c4541 n16__i14__i17__net9 vss 34.6391e-18
c4542 n2__net11 vss 17.2396e-18
c4543 n3__net11 vss 9.69829e-18
c4544 n37__i14__net3 vss 46.7225e-18
c4545 n39__i14__net3 vss 45.9179e-18
c4546 n41__i14__net3 vss 45.3028e-18
c4547 n42__i14__net3 vss 46.4399e-18
c4548 n43__i14__net3 vss 46.7225e-18
c4549 n45__i14__net3 vss 45.012e-18
c4550 n47__i14__net3 vss 44.8034e-18
c4551 n2__y_out_2 vss 9.24549e-18
c4552 n7__x_out_0 vss 9.25955e-18
c4553 n26__i14__i17__net8 vss 103.076e-18
c4554 n16__i14__i17__net11 vss 98.8613e-18
c4555 n17__i14__i17__net11 vss 142.766e-18
c4556 n2__net9 vss 16.6976e-18
c4557 n3__net9 vss 13.717e-18
c4558 n4__net9 vss 17.0059e-18
c4559 n7__i14__i11__net2 vss 90.7819e-18
c4560 n8__i14__i11__net2 vss 63.7124e-18
c4561 n7__i14__i14__net2 vss 91.208e-18
c4562 n8__i14__i14__net2 vss 63.6238e-18
c4563 n7__i14__i15__net2 vss 90.8291e-18
c4564 n8__i14__i15__net2 vss 63.9323e-18
c4565 n7__i14__i12__net2 vss 91.2463e-18
c4566 n8__i14__i12__net2 vss 62.6475e-18
c4567 n658__r_out vss 101.93e-18
c4568 n657__r_out vss 21.2413e-18
c4569 n7__x_out_3 vss 8.92219e-18
c4570 n7__x_out_1 vss 8.47748e-18
c4571 n23__ck vss 18.6756e-18
c4572 n2__i9__i4__net1 vss 16.3029e-18
c4573 n3__i9__i4__net1 vss 8.60249e-18
c4574 n3__i14__clk_div4_out_b vss 293.088e-18
c4575 n2__net12 vss 18.5603e-18
c4576 n3__net12 vss 10.5033e-18
c4577 n2__y_out_3 vss 9.24035e-18
c4578 n2__y_out_1 vss 9.21802e-18
c4579 n2__net10 vss 19.6274e-18
c4580 n3__net10 vss 15.7216e-18
c4581 n4__net10 vss 18.1488e-18
c4582 n7__i14__x_out_b_1 vss 45.2632e-18
c4583 n7__i14__y_out_b_2 vss 44.416e-18
c4584 n7__i14__y_out_b_1 vss 42.91e-18
c4585 n7__i14__x_out_b_0 vss 42.638e-18
c4586 n2__i13__a3 vss 30.4653e-18
c4587 n2__i13__a1 vss 30.4297e-18
c4588 n27__ck vss 12.3297e-18
c4589 n2__i13__a2 vss 25.3455e-18
c4590 n2__i13__a0 vss 25.42e-18
c4591 n52__reset vss 17.1795e-18
c4592 n2__i9__i4__net5 vss 20.0342e-18
c4593 n3__i9__i4__net5 vss 10.256e-18
c4594 n2__i13__i17__net1 vss 11.8495e-18
c4595 n2__i13__i16__net1 vss 11.8509e-18
c4596 n56__reset vss 13.1304e-18
c4597 n5__ck_buff vss 55.7167e-18
c4598 n6__ck_buff vss 36.5908e-18
c4599 n13__ck_b vss 38.8313e-18
c4600 n4__net13 vss 9.57882e-18
c4601 n6__net13 vss 9.26733e-18
c4602 n2__i9__net2 vss 9.80739e-18
c4603 n6__i13__a2 vss 10.7872e-18
c4604 n6__i13__a0 vss 10.728e-18
c4605 n17__y_out_2 vss 43.04e-18
c4606 n17__x_out_0 vss 41.0053e-18
c4607 n8__i13__i14__net2 vss 38.4798e-18
c4608 n9__i13__i14__net2 vss 33.3547e-18
c4609 n7__i13__i12__net2 vss 29.7565e-18
c4610 n11__i13__i12__net2 vss 38.0753e-18
c4611 n12__i13__i14__net2 vss 26.198e-18
c4612 n12__i13__i12__net2 vss 28.4473e-18
c4613 n4__net14 vss 12.0257e-18
c4614 n6__net14 vss 11.5965e-18
c4615 n14__net11 vss 47.5873e-18
c4616 n15__net11 vss 38.0555e-18
c4617 n2__i9__net1 vss 17.7652e-18
c4618 n6__i13__a3 vss 9.4379e-18
c4619 n6__i13__a1 vss 9.17945e-18
c4620 n11__ck4 vss 14.1136e-18
c4621 n4__reset_buff vss 44.5121e-18
c4622 n5__reset_buff vss 45.787e-18
c4623 n12__net9 vss 52.9959e-18
c4624 n2__shift vss 17.5831e-18
c4625 n6__shift vss 14.9646e-18
c4626 n10__shift vss 16.4499e-18
c4627 n2__i13__net11 vss 30.8649e-18
c4628 n2__i13__net12 vss 31.0375e-18
c4629 n7__i9__i4__net2 vss 90.7415e-18
c4630 n8__i9__i4__net2 vss 59.0655e-18
c4631 n2__i13__net1 vss 25.2776e-18
c4632 n2__i13__net2 vss 25.3312e-18
c4633 n16__y_out_3 vss 46.8091e-18
c4634 n17__y_out_1 vss 46.9489e-18
c4635 n8__i13__i15__net2 vss 38.2272e-18
c4636 n9__i13__i15__net2 vss 32.053e-18
c4637 n7__i13__i13__net2 vss 30.2066e-18
c4638 n11__i13__i13__net2 vss 37.8806e-18
c4639 n12__i13__i15__net2 vss 24.5033e-18
c4640 n12__i13__i13__net2 vss 34.9352e-18
c4641 n2__i13__i19__net1 vss 11.5494e-18
c4642 n2__i13__i18__net1 vss 11.5508e-18
c4643 n14__net12 vss 40.8571e-18
c4644 n15__net12 vss 35.332e-18
c4645 n6__i13__net1 vss 10.3899e-18
c4646 n6__i13__net2 vss 10.3307e-18
c4647 n2__i2__net1 vss 10.9335e-18
c4648 n2__i1__net1 vss 10.5797e-18
c4649 n2__i0__net1 vss 10.8867e-18
c4650 n12__net10 vss 42.7989e-18
c4651 n9__i13__i17__net1 vss 57.4577e-18
c4652 n9__i13__i16__net1 vss 57.446e-18
c4653 n12__net13 vss 40.5085e-18
c4654 n6__i13__net11 vss 9.18114e-18
c4655 n6__i13__net12 vss 10.4106e-18
c4656 n5__i9__net2 vss 43.1898e-18
c4657 n12__net14 vss 39.8638e-18
c4658 n2__i13__net7 vss 31.0723e-18
c4659 n2__i13__net17 vss 28.1013e-18
c4660 n23__i13__a3 vss 136.794e-18
c4661 n23__i13__a1 vss 136.194e-18
c4662 n2__i13__net18 vss 25.2229e-18
c4663 n2__i13__net23 vss 23.4708e-18
c4664 n8__i13__i17__i4__net2 vss 38.206e-18
c4665 n9__i13__i17__i4__net2 vss 30.9726e-18
c4666 n7__i13__i16__i4__net2 vss 30.6554e-18
c4667 n11__i13__i16__i4__net2 vss 38.0813e-18
c4668 n12__i13__i17__i4__net2 vss 53.9035e-18
c4669 n12__i13__i16__i4__net2 vss 59.731e-18
c4670 n2__i13__i20__net1 vss 11.3747e-18
c4671 n2__i2__net74 vss 17.1616e-18
c4672 n3__i2__net74 vss 8.90488e-18
c4673 n2__i1__net74 vss 16.4071e-18
c4674 n3__i1__net74 vss 8.62607e-18
c4675 n2__i0__net74 vss 15.9887e-18
c4676 n3__i0__net74 vss 7.87369e-18
c4677 n6__i13__net18 vss 10.2316e-18
c4678 n42__shift vss 77.1891e-18
c4679 n43__shift vss 83.2654e-18
c4680 n44__shift vss 148.502e-18
c4681 n9__i13__i19__net1 vss 56.3092e-18
c4682 n9__i13__i18__net1 vss 59.0097e-18
c4683 n6__i13__net7 vss 11.0916e-18
c4684 n542__vddio vss 88.9792e-18
c4685 n544__vddio vss 64.2755e-18
c4686 n545__vddio vss 78.7853e-18
c4687 n546__vddio vss 78.7853e-18
c4688 n547__vddio vss 62.6718e-18
c4689 n549__vddio vss 69.6614e-18
c4690 n550__vddio vss 78.7853e-18
c4691 n551__vddio vss 69.9514e-18
c4692 n552__vddio vss 53.9195e-18
c4693 n554__vddio vss 69.6614e-18
c4694 n555__vddio vss 78.7853e-18
c4695 n556__vddio vss 78.7492e-18
c4696 n557__vddio vss 62.6718e-18
c4697 n559__vddio vss 93.3856e-18
c4698 n588__vddio vss 69.0565e-18
c4699 n589__vddio vss 69.0565e-18
c4700 n616__vddio vss 126.503e-18
c4701 n619__vddio vss 126.503e-18
c4702 n621__vddio vss 131.491e-18
c4703 n623__vddio vss 131.494e-18
c4704 n628__vddio vss 15.0545e-18
c4705 n2__i2__net76 vss 20.3275e-18
c4706 n3__i2__net76 vss 10.4777e-18
c4707 n2__i1__net76 vss 19.6074e-18
c4708 n3__i1__net76 vss 10.0003e-18
c4709 n2__i0__net76 vss 17.3354e-18
c4710 n3__i0__net76 vss 8.64307e-18
c4711 n19__i13__net11 vss 142.179e-18
c4712 n23__i13__net12 vss 139.872e-18
c4713 n9__i13__i19__i4__net2 vss 32.642e-18
c4714 n12__i13__i19__i4__net2 vss 54.6832e-18
c4715 n12__i13__i18__i4__net2 vss 59.6532e-18
c4716 n2__i2__net73 vss 109.471e-18
c4717 n3__i2__net73 vss 69.7711e-18
c4718 n2__i1__net73 vss 108.076e-18
c4719 n3__i1__net73 vss 69.9024e-18
c4720 n2__i0__net73 vss 110.018e-18
c4721 n3__i0__net73 vss 69.521e-18
c4722 n697__i18__net5 vss 152.08e-18
c4723 n8__serial_out vss 9.8175e-18
c4724 n9__net4 vss 9.53395e-18
c4725 n7__net3 vss 10.1598e-18
c4726 n3__i18__net2 vss 37.5516e-18
c4727 n4__i18__net2 vss 37.5473e-18
c4728 n5__i18__net2 vss 43.3903e-18
c4729 n34__reset_buff vss 47.0768e-18
c4730 n38__reset_buff vss 46.0183e-18
c4731 n9__i13__i20__net1 vss 57.097e-18
c4732 n8__i13__net3 vss 45.2539e-18
c4733 n11__r0 vss 15.1934e-18
c4734 n6__r2 vss 15.1934e-18
c4735 n2__r1 vss 15.1934e-18
c4736 n3__i18__net1 vss 42.9807e-18
c4737 n7__i2__net75 vss 91.6704e-18
c4738 n8__i2__net75 vss 56.1793e-18
c4739 n7__i1__net75 vss 90.1123e-18
c4740 n8__i1__net75 vss 55.2002e-18
c4741 n7__i0__net75 vss 91.1685e-18
c4742 n8__i0__net75 vss 61.4249e-18
c4743 n19__i13__net7 vss 147.061e-18
c4744 n2__net7 vss 17.4798e-18
c4745 n3__net7 vss 17.7691e-18
c4746 n4__net7 vss 9.83273e-18
c4747 n2__net6 vss 17.118e-18
c4748 n3__net6 vss 17.4354e-18
c4749 n4__net6 vss 10.3289e-18
c4750 n2__net8 vss 15.9146e-18
c4751 n3__net8 vss 13.9478e-18
c4752 n4__net8 vss 9.38016e-18
c4753 n8__i13__i20__i4__net2 vss 38.0644e-18
c4754 n9__i13__i20__i4__net2 vss 32.0293e-18
c4755 n12__i13__i20__i4__net2 vss 57.346e-18
c4756 n207__i18__net4 vss 133.978e-18
c4757 n640__vddio vss 10.22e-18
c4758 n641__vddio vss 15.3233e-18
c4759 n649__vddio vss 19.2765e-18
c4760 n9__serial_out_b_high vss 121.666e-18
c4761 n20__serial_out vss 42.9279e-18
c4762 n12__net4 vss 43.1531e-18
c4763 n10__net3 vss 42.5787e-18
c4764 n53__i18__net3 vss 57.9768e-18
c4765 n54__i18__net3 vss 103.325e-18
c4766 n6__i12__bio vss 98.7306e-18
c4767 n14__i18__net2 vss 76.0474e-18
c4768 n12__i12__bcore_bar vss 96.5209e-18
c4769 n34__vdd vss 53.3644e-18
c4770 n35__vdd vss 65.566e-18
c4771 n36__vdd vss 53.2166e-18
c4772 n37__vdd vss 33.9098e-18
c4773 n39__vdd vss 166.738e-18
c4774 n41__vdd vss 140.164e-18
c4775 n43__vdd vss 32.3532e-18
c4776 n44__vdd vss 55.8261e-18
c4777 n45__vdd vss 106.676e-18
c4778 n47__vdd vss 180.21e-18
c4779 n49__vdd vss 109.878e-18
c4780 n50__vdd vss 76.4966e-18
c4781 n51__vdd vss 34.1195e-18
c4782 n53__vdd vss 32.4429e-18
c4783 n54__vdd vss 49.9589e-18
c4784 n55__vdd vss 39.0007e-18
c4785 n56__vdd vss 110.202e-18
c4786 n58__vdd vss 28.3578e-18
c4787 n59__vdd vss 88.9536e-18
c4788 n60__vdd vss 177.546e-18
c4789 n62__vdd vss 64.1675e-18
c4790 n63__vdd vss 37.1824e-18
c4791 n64__vdd vss 27.8857e-18
c4792 n65__vdd vss 44.1276e-18
c4793 n66__vdd vss 30.6493e-18
c4794 n118__vdd vss 74.1071e-18
c4795 n121__vdd vss 55.0296e-18
c4796 n125__vdd vss 274.621e-18
c4797 n11__net7 vss 40.9021e-18
c4798 n11__net6 vss 43.3554e-18
c4799 n11__net8 vss 41.1244e-18
c4800 n671__vddio vss 33.108e-18
c4801 n674__vddio vss 96.6579e-18
c4802 n8__i18__net1 vss 75.0791e-18
c4803 n9__r0_buff vss 41.6847e-18
c4804 n10__r0_buff vss 50.0139e-18
c4805 n9__r2_buff vss 38.1819e-18
c4806 n13__r2_buff vss 48.3021e-18
c4807 n9__r1_buff vss 41.3763e-18
c4808 n10__r1_buff vss 46.6962e-18
c4809 n136__vdd vss 37.5121e-18
c4810 n138__vdd vss 22.2929e-18
c4811 n139__vdd vss 27.5674e-18
c4812 n141__vdd vss 8.33144e-18
c4813 n142__vdd vss 15.5043e-18
c4814 n143__vdd vss 23.7985e-18
c4815 n144__vdd vss 18.359e-18
c4816 n146__vdd vss 76.0906e-18
c4817 n147__vdd vss 65.8013e-18
c4818 n148__vdd vss 32.9553e-18
c4819 n150__vdd vss 149.05e-18
c4820 n151__vdd vss 138.374e-18
c4821 n152__vdd vss 124.346e-18
c4822 n153__vdd vss 21.9475e-18
c4823 n154__vdd vss 18.9017e-18
c4824 n156__vdd vss 37.0805e-18
c4825 n157__vdd vss 53.7294e-18
c4826 n158__vdd vss 7.35168e-18
c4827 n161__vdd vss 54.2775e-18
c4828 n162__vdd vss 26.2182e-18
c4829 n164__vdd vss 58.9566e-18
c4830 n165__vdd vss 30.4118e-18
c4831 n166__vdd vss 33.3863e-18
c4832 n168__vdd vss 35.8801e-18
c4833 n169__vdd vss 29.0505e-18
c4834 n170__vdd vss 37.8701e-18
c4835 n171__vdd vss 30.9927e-18
c4836 n173__vdd vss 23.8404e-18
c4837 n174__vdd vss 70.2996e-18
c4838 n175__vdd vss 31.7414e-18
c4839 n177__vdd vss 63.6026e-18
c4840 n178__vdd vss 47.3763e-18
c4841 n179__vdd vss 51.1469e-18
c4842 n181__vdd vss 26.4741e-18
c4843 n182__vdd vss 36.3632e-18
c4844 n183__vdd vss 22.5198e-18
c4845 n184__vdd vss 39.7463e-18
c4846 n186__vdd vss 90.2831e-18
c4847 n187__vdd vss 29.3237e-18
c4848 n189__vdd vss 52.0073e-18
c4849 n190__vdd vss 60.5455e-18
c4850 n191__vdd vss 48.6829e-18
c4851 n192__vdd vss 59.1246e-18
c4852 n193__vdd vss 26.756e-18
c4853 n195__vdd vss 86.2875e-18
c4854 n196__vdd vss 74.1156e-18
c4855 n198__vdd vss 23.5787e-18
c4856 n199__vdd vss 43.0661e-18
c4857 n200__vdd vss 32.0266e-18
c4858 n201__vdd vss 57.5462e-18
c4859 n202__vdd vss 39.6558e-18
c4860 n203__vdd vss 64.8731e-18
c4861 n205__vdd vss 36.1786e-18
c4862 n206__vdd vss 87.065e-18
c4863 n207__vdd vss 147.863e-18
c4864 n209__vdd vss 115.17e-18
c4865 n292__vdd vss 34.2149e-18
c4866 n295__vdd vss 41.9353e-18
c4867 n297__vdd vss 59.7855e-18
c4868 n298__vdd vss 70.1506e-18
c4869 n300__vdd vss 12.6776e-18
c4870 n301__vdd vss 32.5817e-18
c4871 n302__vdd vss 50.6922e-18
c4872 n303__vdd vss 31.1928e-18
c4873 n305__vdd vss 171.027e-18
c4874 n306__vdd vss 156.276e-18
c4875 n307__vdd vss 76.6108e-18
c4876 n309__vdd vss 338.757e-18
c4877 n310__vdd vss 457.906e-18
c4878 n311__vdd vss 218.784e-18
c4879 n312__vdd vss 50.6163e-18
c4880 n314__vdd vss 25.3528e-18
c4881 n316__vdd vss 22.1875e-18
c4882 n317__vdd vss 10.1163e-18
c4883 n319__vdd vss 3.18074e-18
c4884 n321__vdd vss 13.9421e-18
c4885 n322__vdd vss 7.11357e-18
c4886 n324__vdd vss 80.0874e-18
c4887 n325__vdd vss 87.1179e-18
c4888 n326__vdd vss 35.0032e-18
c4889 n328__vdd vss 32.4506e-18
c4890 n329__vdd vss 49.9589e-18
c4891 n330__vdd vss 39.3429e-18
c4892 n331__vdd vss 110.224e-18
c4893 n333__vdd vss 28.3517e-18
c4894 n334__vdd vss 89.0033e-18
c4895 n335__vdd vss 177.413e-18
c4896 n337__vdd vss 64.2022e-18
c4897 n338__vdd vss 36.6396e-18
c4898 n339__vdd vss 28.1729e-18
c4899 n340__vdd vss 44.1245e-18
c4900 n341__vdd vss 30.6306e-18
c4901 n343__vdd vss 54.8774e-18
c4902 n344__vdd vss 99.8044e-18
c4903 n345__vdd vss 54.9721e-18
c4904 n347__vdd vss 274.671e-18
c4905 n679__vddio vss 56.2611e-18
c4906 n698__vddio vss 20.5587e-18
c4907 n701__vddio vss 39.1762e-18
c4908 n702__vddio vss 39.6935e-18
c4909 n703__vddio vss 25.3107e-18
c4910 n705__vddio vss 33.6018e-18
c4911 n706__vddio vss 39.6935e-18
c4912 n707__vddio vss 30.1815e-18
c4913 n709__vddio vss 25.2556e-18
c4914 n710__vddio vss 39.6935e-18
c4915 n711__vddio vss 39.6935e-18
c4916 n713__vddio vss 38.2337e-18
c4917 n714__vddio vss 39.6935e-18
c4918 n715__vddio vss 27.5486e-18
c4919 n717__vddio vss 28.3361e-18
c4920 n718__vddio vss 39.6935e-18
c4921 n719__vddio vss 35.9475e-18
c4922 n721__vddio vss 43.4945e-18
c4923 n722__vddio vss 39.6935e-18
c4924 n723__vddio vss 39.6935e-18
c4925 n724__vddio vss 25.3107e-18
c4926 n726__vddio vss 30.9689e-18
c4927 n727__vddio vss 39.6935e-18
c4928 n728__vddio vss 32.8144e-18
c4929 n730__vddio vss 25.2556e-18
c4930 n731__vddio vss 39.6935e-18
c4931 n732__vddio vss 39.6935e-18
c4932 n733__vddio vss 25.3107e-18
c4933 n735__vddio vss 33.6018e-18
c4934 n736__vddio vss 39.6935e-18
c4935 n737__vddio vss 30.1815e-18
c4936 n739__vddio vss 25.2556e-18
c4937 n740__vddio vss 39.6935e-18
c4938 n741__vddio vss 39.6935e-18
c4939 n743__vddio vss 38.2337e-18
c4940 n744__vddio vss 39.6935e-18
c4941 n745__vddio vss 27.5486e-18
c4942 n747__vddio vss 28.3361e-18
c4943 n748__vddio vss 39.6935e-18
c4944 n749__vddio vss 35.9475e-18
c4945 n751__vddio vss 43.4945e-18
c4946 n752__vddio vss 39.6935e-18
c4947 n753__vddio vss 39.6935e-18
c4948 n754__vddio vss 25.3107e-18
c4949 n756__vddio vss 30.9689e-18
c4950 n757__vddio vss 39.6935e-18
c4951 n758__vddio vss 32.8144e-18
c4952 n760__vddio vss 25.2556e-18
c4953 n761__vddio vss 53.9446e-18
c4954 n964__vddio vss 8.3925e-18
rc1 r_out n458__r_out 4.822e-3
rc2 vddio n1022__vddio 460.5e-3
rc3 n1022__vddio n1021__vddio 227.4e-3
rc5 n1021__vddio n1024__vddio 3.418e-3
rc6 n1024__vddio vddio 4.656e-3
rc7 vddio n1025__vddio 5.445e-3
rc8 n1025__vddio n1012__vddio 53.55e-3
rc9 n439__vddio n1022__vddio 46.67e-3
rc10 n1015__vddio n1021__vddio 46.67e-3
rc11 n1014__vddio n1024__vddio 46.67e-3
rc12 n1013__vddio n1025__vddio 46.67e-3
rc13 vdd n30__vdd 90.94e-3
rc14 n30__vdd n19__vdd 244.6e-3
rc15 n19__vdd vdd 371e-3
rc16 n1342__vss n1343__vss 2.725e-3
rc17 n1343__vss vss 4.921e-3
rc19 vss n1345__vss 4.723e-3
rc20 n1345__vss n622__vss 150.5e-3
rc21 n622__vss n464__vss 90.82e-3
rc22 n464__vss n457__vss 22.03e-3
rc23 n457__vss vss 435.9e-3
rc24 vss n1346__vss 437.5e-3
rc25 n1346__vss n1347__vss 22.03e-3
rc26 n1347__vss n1348__vss 90.82e-3
rc27 n1348__vss n1349__vss 67.12e-3
rc28 n1349__vss n1342__vss 146.9e-3
rc29 n1334__vss n1342__vss 46.67e-3
rc30 n1335__vss n1343__vss 46.67e-3
rc31 n1336__vss vss 46.67e-3
rc32 n1337__vss n1345__vss 46.67e-3
rc33 n456__vss n1346__vss 46.67e-3
rc34 n459__vss n1347__vss 46.67e-3
rc35 n621__vss n1348__vss 46.67e-3
rd1 n458__r_out n459__r_out 65e-3
rd2 n14__vdd n19__vdd 73.44e-3
rd3 n14__vdd n15__vdd 121.2e-3
rd4 n15__vdd n18__vdd 121.2e-3
rd5 n452__vss n453__vss 204.5e-3
rd6 n453__vss n454__vss 121.2e-3
rd7 n454__vss n455__vss 121.2e-3
rd8 n455__vss n456__vss 33.83e-3
rd9 n456__vss n457__vss 226.6e-3
rd10 n435__vddio n436__vddio 170.1e-3
rd11 n436__vddio n437__vddio 77e-3
rd12 n437__vddio n438__vddio 42.96e-3
rd13 n438__vddio n439__vddio 33e-3
rd14 n439__vddio n440__vddio 83.33e-3
rd15 n458__vss n459__vss 109.3e-3
rd17 n459__vss n461__vss 34.24e-3
rd18 n461__vss n462__vss 61.85e-3
rd19 n462__vss n463__vss 61.43e-3
rd20 n463__vss n464__vss 76.55e-3
rd21 n619__vss n620__vss 137.3e-3
rd22 n620__vss n621__vss 38.21e-3
rd23 n621__vss n622__vss 251.7e-3
rd24 n30__vdd n29__vdd 367.7e-3
rd25 n1010__vddio n1011__vddio 188.2e-3
rd26 n1011__vddio n1012__vddio 314.6e-3
rd28 n1012__vddio n1013__vddio 86.54e-3
rd30 n1013__vddio n1014__vddio 77e-3
rd32 n1014__vddio n1015__vddio 42.96e-3
rd34 n1015__vddio n1016__vddio 33e-3
rd35 n1016__vddio n1021__vddio 46.67e-3
rd36 n1333__vss n1334__vss 25.94e-3
rd38 n1334__vss n1335__vss 34.24e-3
rd40 n1335__vss n1336__vss 61.85e-3
rd42 n1336__vss n1337__vss 61.43e-3
re2 n13__vdd n14__vdd 166.7e-3
re3 n15__vdd n16__vdd 166.7e-3
re4 n17__vdd n18__vdd 166.7e-3
re5 n425__vss n452__vss 83.33e-3
re6 n453__vss n426__vss 166.7e-3
re7 n427__vss n454__vss 166.7e-3
re8 n455__vss n428__vss 166.7e-3
re9 n435__vddio n441__vddio 83.33e-3
re10 n442__vddio n436__vddio 166.7e-3
re11 n437__vddio n443__vddio 166.7e-3
re12 n444__vddio n438__vddio 166.7e-3
re13 n440__vddio n445__vddio 83.33e-3
re14 n465__vss n458__vss 83.33e-3
re15 n459__vss n466__vss 166.7e-3
re16 n467__vss n461__vss 166.7e-3
re17 n462__vss n468__vss 166.7e-3
re18 n469__vss n463__vss 166.7e-3
re19 n617__vss n619__vss 83.33e-3
re20 n620__vss n618__vss 83.33e-3
re21 n29__vdd n28__vdd 83.33e-3
re22 n427__vdd n428__vdd 390.1e-3
re23 n1003__vddio n1010__vddio 83.33e-3
re24 n1011__vddio n1004__vddio 83.33e-3
re25 n1005__vddio n1012__vddio 83.33e-3
re26 n1013__vddio n1006__vddio 83.33e-3
re27 n1007__vddio n1014__vddio 83.33e-3
re28 n1015__vddio n1008__vddio 83.33e-3
re29 n1009__vddio n1016__vddio 83.33e-3
re30 n1333__vss n1328__vss 83.33e-3
re31 n1329__vss n1334__vss 83.33e-3
re32 n1335__vss n1330__vss 83.33e-3
re33 n1331__vss n1336__vss 83.33e-3
re34 n1337__vss n1332__vss 83.33e-3
rf1 n459__r_out n430__r_out 41.67e-3
rf2 n10__vdd n13__vdd 83.33e-3
rf3 n16__vdd n11__vdd 83.33e-3
rf4 n12__vdd n17__vdd 83.33e-3
rf19 n615__vss n617__vss 83.33e-3
rf20 n618__vss n616__vss 83.33e-3
rf21 n28__vdd n27__vdd 83.33e-3
rf22 n427__vdd n425__vdd 83.33e-3
rf23 n426__vdd n428__vdd 83.33e-3
rf24 n996__vddio n1003__vddio 83.33e-3
rf25 n1004__vddio n997__vddio 83.33e-3
rf26 n998__vddio n1005__vddio 83.33e-3
rf27 n1006__vddio n999__vddio 83.33e-3
rf28 n1000__vddio n1007__vddio 83.33e-3
rf29 n1008__vddio n1001__vddio 83.33e-3
rf30 n1002__vddio n1009__vddio 83.33e-3
rf31 n1328__vss n1323__vss 83.33e-3
rf32 n1324__vss n1329__vss 83.33e-3
rf33 n1330__vss n1325__vss 83.33e-3
rf34 n1326__vss n1331__vss 83.33e-3
rf35 n1332__vss n1327__vss 83.33e-3
rg1 n430__r_out n431__r_out 83.33e-3
rg5 n413__vss n425__vss 83.33e-3
rg6 n426__vss n414__vss 83.33e-3
rg7 n415__vss n427__vss 83.33e-3
rg8 n428__vss n416__vss 83.33e-3
rg9 n441__vddio n421__vddio 83.33e-3
rg10 n422__vddio n442__vddio 83.33e-3
rg11 n443__vddio n425__vddio 83.33e-3
rg12 n426__vddio n444__vddio 83.33e-3
rg13 n445__vddio n428__vddio 83.33e-3
rg14 n440__vss n465__vss 83.33e-3
rg15 n466__vss n442__vss 83.33e-3
rg16 n443__vss n467__vss 83.33e-3
rg17 n468__vss n446__vss 83.33e-3
rg18 n447__vss n469__vss 83.33e-3
rg19 n59__reset n50__reset 1.9998
rg20 n615__vss n509__vss 83.33e-3
rg21 n510__vss n616__vss 83.33e-3
rg22 n37__ck n33__ck 427.7e-3
rg23 n33__ck n20__ck 6.0231
rg24 ck n37__ck 19.99e-3
rg27 reset n66__reset 1.3364
rg28 n26__vdd n27__vdd 83.33e-3
rg29 n423__vdd n425__vdd 83.33e-3
rg30 n426__vdd n424__vdd 83.33e-3
rg31 n996__vddio n989__vddio 83.33e-3
rg32 n990__vddio n997__vddio 83.33e-3
rg33 n998__vddio n991__vddio 83.33e-3
rg34 n992__vddio n999__vddio 83.33e-3
rg35 n1000__vddio n993__vddio 83.33e-3
rg36 n994__vddio n1001__vddio 83.33e-3
rg37 n1002__vddio n995__vddio 83.33e-3
rg38 n1318__vss n1323__vss 83.33e-3
rg39 n1324__vss n1319__vss 83.33e-3
rg40 n1320__vss n1325__vss 83.33e-3
rg41 n1326__vss n1321__vss 83.33e-3
rg42 n1322__vss n1327__vss 83.33e-3
rh1 x3 n5__x3 39.86e-3
rh2 x2 n5__x2 39.86e-3
rh3 x1 n5__x1 39.86e-3
rh4 x0 n5__x0 39.86e-3
rh5 n19__ck n20__ck 500e-3
rh6 n7__vdd n10__vdd 83.33e-3
rh7 n11__vdd n8__vdd 83.33e-3
rh8 n9__vdd n12__vdd 83.33e-3
rh9 n14__i14__i17__net7 n9__i14__i17__net7 1.7125
rh10 n22__i14__i17__net1 n12__i14__i17__net1 2.6048
rh11 n25__i14__i17__net1 n21__i14__i17__net1 249.3e-3
rh12 n4__y3 y3 2.8864
rh13 n5__y2 y2 2.8804
rh14 n4__y1 y1 2.8804
rh15 n5__y0 y0 2.8297
rh16 n16__i14__i17__net7 n13__i14__i17__net7 646.6e-3
rh17 n47__reset n13__reset 3.4599
rh18 n413__vss n409__vss 83.33e-3
rh19 n410__vss n414__vss 83.33e-3
rh20 n415__vss n411__vss 83.33e-3
rh21 n412__vss n416__vss 83.33e-3
rh22 n654__r_out n641__r_out 127.5e-3
rh23 n641__r_out n628__r_out 125.7e-3
rh24 n628__r_out n615__r_out 126.6e-3
rh25 n615__r_out n602__r_out 127.5e-3
rh26 n602__r_out n587__r_out 124.8e-3
rh27 n587__r_out n576__r_out 127.5e-3
rh28 n576__r_out n563__r_out 125.7e-3
rh29 n563__r_out n550__r_out 126.6e-3
rh30 n550__r_out n537__r_out 127.5e-3
rh31 n537__r_out n524__r_out 126.6e-3
rh32 n524__r_out n504__r_out 127.5e-3
rh33 n504__r_out n491__r_out 125.7e-3
rh34 n491__r_out n485__r_out 126.6e-3
rh35 n485__r_out n472__r_out 127.5e-3
rh36 n472__r_out n456__r_out 126.6e-3
rh37 n456__r_out n436__r_out 127.5e-3
rh38 n436__r_out n428__r_out 125.7e-3
rh39 n428__r_out n415__r_out 126.6e-3
rh40 n415__r_out n402__r_out 127.5e-3
rh41 n402__r_out n389__r_out 124.8e-3
rh42 n389__r_out n369__r_out 127.5e-3
rh43 n369__r_out n363__r_out 125.7e-3
rh44 n363__r_out n350__r_out 126.6e-3
rh45 n350__r_out n330__r_out 127.5e-3
rh46 n330__r_out n317__r_out 126.6e-3
rh47 n317__r_out n304__r_out 127.5e-3
rh48 n304__r_out n291__r_out 125.7e-3
rh49 n291__r_out n285__r_out 126.6e-3
rh50 n285__r_out n265__r_out 127.5e-3
rh51 n265__r_out n252__r_out 125.7e-3
rh52 n252__r_out n239__r_out 127.5e-3
rh53 n239__r_out n226__r_out 125.7e-3
rh54 n226__r_out n220__r_out 126.6e-3
rh55 n220__r_out n200__r_out 127.5e-3
rh56 n200__r_out n194__r_out 124.8e-3
rh57 n194__r_out n656__r_out 42.03e-3
rh58 n656__r_out n431__r_out 597.5e-3
rh59 n431__r_out n657__r_out 69.03e-3
rh60 n657__r_out n175__r_out 86.69e-3
rh61 n175__r_out n169__r_out 133.3e-3
rh62 n169__r_out n156__r_out 134.2e-3
rh63 n156__r_out n143__r_out 135.2e-3
rh64 n143__r_out n123__r_out 134.2e-3
rh65 n123__r_out n110__r_out 135.2e-3
rh66 n110__r_out n97__r_out 133.3e-3
rh67 n97__r_out n91__r_out 134.2e-3
rh68 n91__r_out n71__r_out 135.2e-3
rh69 n71__r_out n65__r_out 132.3e-3
rh70 n65__r_out n45__r_out 135.2e-3
rh71 n45__r_out n39__r_out 133.3e-3
rh72 n39__r_out n26__r_out 134.2e-3
rh73 n26__r_out n6__r_out 135.2e-3
rh74 n657__r_out n195__r_out 44.51e-3
rh75 n195__r_out n201__r_out 132.3e-3
rh76 n201__r_out n221__r_out 135.2e-3
rh77 n221__r_out n227__r_out 134.2e-3
rh78 n227__r_out n240__r_out 133.3e-3
rh79 n240__r_out n253__r_out 135.2e-3
rh80 n253__r_out n266__r_out 133.3e-3
rh81 n266__r_out n286__r_out 135.2e-3
rh82 n286__r_out n292__r_out 134.2e-3
rh83 n292__r_out n305__r_out 133.3e-3
rh84 n305__r_out n318__r_out 135.2e-3
rh85 n318__r_out n331__r_out 134.2e-3
rh86 n331__r_out n351__r_out 135.2e-3
rh87 n351__r_out n364__r_out 134.2e-3
rh88 n364__r_out n370__r_out 133.3e-3
rh89 n370__r_out n390__r_out 135.2e-3
rh90 n390__r_out n403__r_out 132.3e-3
rh91 n403__r_out n416__r_out 135.2e-3
rh92 n416__r_out n429__r_out 134.2e-3
rh93 n429__r_out n437__r_out 133.3e-3
rh94 n437__r_out n457__r_out 135.2e-3
rh95 n457__r_out n473__r_out 134.2e-3
rh96 n473__r_out n486__r_out 135.2e-3
rh97 n486__r_out n492__r_out 134.2e-3
rh98 n492__r_out n505__r_out 133.3e-3
rh99 n505__r_out n525__r_out 135.2e-3
rh100 n525__r_out n538__r_out 134.2e-3
rh101 n538__r_out n551__r_out 135.2e-3
rh102 n551__r_out n564__r_out 134.2e-3
rh103 n564__r_out n577__r_out 133.3e-3
rh104 n577__r_out n590__r_out 135.2e-3
rh105 n590__r_out n603__r_out 132.3e-3
rh106 n603__r_out n616__r_out 135.2e-3
rh107 n616__r_out n629__r_out 134.2e-3
rh108 n629__r_out n642__r_out 133.3e-3
rh109 n642__r_out n655__r_out 135.2e-3
rh110 n6__r_out n5__r_out 772.8e-3
rh111 n5__r_out n25__r_out 127.5e-3
rh112 n25__r_out n38__r_out 126.6e-3
rh113 n38__r_out n44__r_out 125.7e-3
rh114 n44__r_out n64__r_out 127.5e-3
rh115 n64__r_out n70__r_out 124.8e-3
rh116 n70__r_out n90__r_out 127.5e-3
rh117 n90__r_out n96__r_out 126.6e-3
rh118 n96__r_out n109__r_out 125.7e-3
rh119 n109__r_out n122__r_out 127.5e-3
rh120 n122__r_out n142__r_out 126.6e-3
rh121 n142__r_out n155__r_out 127.5e-3
rh122 n155__r_out n168__r_out 126.6e-3
rh123 n168__r_out n174__r_out 125.7e-3
rh124 n174__r_out n658__r_out 34.91e-3
rh125 n658__r_out n656__r_out 46.92e-3
rh126 n62__i14__net4 n9__i14__net4 3.4163
rh127 n64__i14__net4 n12__i14__net4 3.4163
rh128 n66__i14__net4 n13__i14__net4 3.4163
rh129 n68__i14__net4 n16__i14__net4 3.4163
rh130 n64__i14__net3 n53__i14__net3 1.5906
rh131 n53__i14__net3 n17__i14__net3 3.3499
rh132 n65__i14__net3 n54__i14__net3 1.5906
rh133 n54__i14__net3 n18__i14__net3 3.3499
rh134 n66__i14__net3 n55__i14__net3 1.5906
rh135 n55__i14__net3 n19__i14__net3 3.3499
rh136 n67__i14__net3 n56__i14__net3 1.0906
rh137 n56__i14__net3 n20__i14__net3 3.3499
rh138 n413__vddio n421__vddio 166.7e-3
rh139 n422__vddio n414__vddio 166.7e-3
rh140 n415__vddio n425__vddio 166.7e-3
rh141 n426__vddio n416__vddio 166.7e-3
rh142 n419__vddio n428__vddio 83.33e-3
rh143 n440__vss n439__vss 83.33e-3
rh144 n435__vss n442__vss 166.7e-3
rh145 n443__vss n436__vss 166.7e-3
rh146 n437__vss n446__vss 166.7e-3
rh147 n447__vss n438__vss 166.7e-3
rh148 n82__i14__net9 n69__i14__net9 2.261
rh149 n69__i14__net9 n29__i14__net9 3.163
rh150 n83__i14__net9 n70__i14__net9 2.261
rh151 n70__i14__net9 n30__i14__net9 3.163
rh152 n84__i14__net9 n71__i14__net9 2.261
rh153 n71__i14__net9 n31__i14__net9 3.163
rh154 n85__i14__net9 n72__i14__net9 1.761
rh155 n72__i14__net9 n32__i14__net9 3.163
rh156 n13__x_out_3 n5__x_out_3 2.3865
rh157 n12__x_out_2 n5__x_out_2 2.3865
rh158 n13__x_out_1 n5__x_out_1 2.3865
rh159 n10__x_out_0 n5__x_out_0 2.3865
rh164 n39__i14__net7 n36__i14__net7 220.1e-3
rh165 n36__i14__net7 n31__i14__net7 781.2e-3
rh166 n38__i14__net11 n35__i14__net11 198.1e-3
rh167 n35__i14__net11 n29__i14__net11 707.9e-3
rh168 n109__i14__net10 n89__i14__net10 3.0271
rh169 n89__i14__net10 n45__i14__net10 2.9799
rh170 n110__i14__net10 n90__i14__net10 3.0271
rh171 n90__i14__net10 n46__i14__net10 2.9799
rh172 n111__i14__net10 n91__i14__net10 3.0271
rh173 n91__i14__net10 n47__i14__net10 2.9799
rh174 n112__i14__net10 n92__i14__net10 2.5271
rh175 n92__i14__net10 n48__i14__net10 2.9799
rh176 n50__reset n25__reset 5.0284
rh177 n13__y_out_0 n8__y_out_0 319.8e-3
rh178 n13__x_out_0 n11__x_out_0 1.0395
rh179 n20__x_out_2 n15__x_out_2 203.2e-3
rh180 n19__x_out_2 n13__x_out_2 1.1454
rh181 n16__y_out_2 n10__y_out_2 196.6e-3
rh182 n15__y_out_2 n6__y_out_2 650.4e-3
rh183 n14__x_out_3 n12__x_out_3 2.0849
rh184 n8__reset_buff n7__reset_buff 217.4e-3
rh185 n10__y_out_3 n5__y_out_3 1.6005
rh186 n32__ck n33__ck 500e-3
rh187 n16__y_out_1 n10__y_out_1 104.1e-3
rh188 n15__y_out_1 n5__y_out_1 1.9474
rh189 n20__x_out_1 n12__x_out_1 2.4901
rh190 n21__x_out_1 n15__x_out_1 306.7e-3
rh191 n21__i13__a2 n19__i13__a2 1.0488
rh192 n22__i13__a0 n20__i13__a0 1.0529
rh193 n509__vss n507__vss 83.33e-3
rh194 n508__vss n510__vss 83.33e-3
rh195 n36__ck n37__ck 250e-3
rh196 n66__reset n59__reset 1.5051
rh197 n62__reset reset 250e-3
rh198 reset n65__reset 250e-3
rh199 n19__reset_buff n9__reset_buff 2.137
rh200 n7__r2_buff r2_buff 744.8e-3
rh201 n7__r1_buff r1_buff 840.9e-3
rh202 n7__r0_buff r0_buff 918.1e-3
rh203 n25__vdd n26__vdd 83.33e-3
rh204 n6__net4 n3__net4 912.2e-3
rh205 n695__i18__net5 n675__i18__net5 127.5e-3
rh206 n675__i18__net5 n669__i18__net5 125.7e-3
rh207 n669__i18__net5 n656__i18__net5 126.6e-3
rh208 n656__i18__net5 n632__i18__net5 127.5e-3
rh209 n632__i18__net5 n630__i18__net5 124.8e-3
rh210 n630__i18__net5 n617__i18__net5 127.5e-3
rh211 n617__i18__net5 n597__i18__net5 125.7e-3
rh212 n597__i18__net5 n591__i18__net5 126.6e-3
rh213 n591__i18__net5 n578__i18__net5 127.5e-3
rh214 n578__i18__net5 n558__i18__net5 126.6e-3
rh215 n558__i18__net5 n552__i18__net5 127.5e-3
rh216 n552__i18__net5 n539__i18__net5 125.7e-3
rh217 n539__i18__net5 n526__i18__net5 126.6e-3
rh218 n526__i18__net5 n513__i18__net5 127.5e-3
rh219 n513__i18__net5 n697__i18__net5 318.7e-3
rh220 n697__i18__net5 n500__i18__net5 396.9e-3
rh221 n697__i18__net5 n514__i18__net5 585.4e-3
rh222 n514__i18__net5 n527__i18__net5 182.9e-3
rh223 n527__i18__net5 n540__i18__net5 181.6e-3
rh224 n540__i18__net5 n553__i18__net5 180.3e-3
rh225 n553__i18__net5 n559__i18__net5 182.9e-3
rh226 n559__i18__net5 n579__i18__net5 181.6e-3
rh227 n579__i18__net5 n592__i18__net5 182.9e-3
rh228 n592__i18__net5 n598__i18__net5 181.6e-3
rh229 n598__i18__net5 n618__i18__net5 180.3e-3
rh230 n618__i18__net5 n631__i18__net5 182.9e-3
rh231 n631__i18__net5 n635__i18__net5 179e-3
rh232 n635__i18__net5 n657__i18__net5 182.9e-3
rh233 n657__i18__net5 n670__i18__net5 181.6e-3
rh234 n670__i18__net5 n676__i18__net5 180.3e-3
rh235 n676__i18__net5 n696__i18__net5 182.9e-3
rh236 n31__ck_b n15__ck_b 4.0005
rh237 n28__reset_buff n16__reset_buff 2.1663
rh238 n37__ck_buff n23__ck_buff 1.7613
rh239 n23__ck_buff n8__ck_buff 2.0622
rh240 n21__reset_b n5__reset_b 4.4405
rh241 n5__reset_b n3__reset_b 242.1e-3
rh242 n205__i18__net4 n194__i18__net4 127.5e-3
rh243 n194__i18__net4 n174__i18__net4 125.7e-3
rh244 n174__i18__net4 n172__i18__net4 126.6e-3
rh245 n172__i18__net4 n161__i18__net4 127.5e-3
rh246 n161__i18__net4 n207__i18__net4 343.8e-3
rh247 n207__i18__net4 n150__i18__net4 318.4e-3
rh248 n207__i18__net4 n162__i18__net4 609.6e-3
rh249 n162__i18__net4 n173__i18__net4 182.9e-3
rh250 n173__i18__net4 n177__i18__net4 181.6e-3
rh251 n177__i18__net4 n195__i18__net4 180.3e-3
rh252 n195__i18__net4 n206__i18__net4 182.9e-3
rh253 n17__net4 n7__net4 3.3813
rh254 n15__net3 n3__net3 3.8713
rh255 n423__vdd n421__vdd 83.33e-3
rh256 n422__vdd n424__vdd 83.33e-3
rh257 n32__serial_out n30__serial_out 459e-3
rh258 n31__serial_out serial_out 463.9e-3
rh259 serial_out n29__serial_out 459e-3
rh260 n17__serial_out_b_high n16__serial_out_b_high 2.067
rh261 n976__vddio n989__vddio 83.33e-3
rh262 n990__vddio n977__vddio 83.33e-3
rh263 n971__vddio n991__vddio 166.7e-3
rh264 n992__vddio n972__vddio 166.7e-3
rh265 n973__vddio n993__vddio 166.7e-3
rh266 n994__vddio n974__vddio 166.7e-3
rh267 n978__vddio n995__vddio 83.33e-3
rh268 n17__r2_buff n2__r2_buff 7.0572
rh269 n16__r1_buff n2__r1_buff 7.0509
rh270 n16__r0_buff n2__r0_buff 8.0627
rh271 n1309__vss n1318__vss 83.33e-3
rh272 n1319__vss n1305__vss 166.7e-3
rh273 n1306__vss n1320__vss 166.7e-3
rh274 n1321__vss n1307__vss 166.7e-3
rh275 n1308__vss n1322__vss 166.7e-3
ri1 n5__r_out n2__r_out 500e-3
ri2 n3__r_out n6__r_out 500e-3
ri3 n25__r_out n23__r_out 500e-3
ri4 n24__r_out n26__r_out 500e-3
ri5 n38__r_out n28__r_out 500e-3
ri6 n29__r_out n39__r_out 500e-3
ri7 n44__r_out n41__r_out 500e-3
ri8 n42__r_out n45__r_out 500e-3
ri9 n64__r_out n54__r_out 500e-3
ri10 n55__r_out n65__r_out 500e-3
ri11 n70__r_out n67__r_out 500e-3
ri12 n68__r_out n71__r_out 500e-3
ri13 n90__r_out n88__r_out 500e-3
ri14 n89__r_out n91__r_out 500e-3
ri15 n96__r_out n93__r_out 500e-3
ri16 n94__r_out n97__r_out 500e-3
ri17 n109__r_out n106__r_out 500e-3
ri18 n107__r_out n110__r_out 500e-3
ri19 n122__r_out n119__r_out 500e-3
ri20 n120__r_out n123__r_out 500e-3
ri21 n142__r_out n140__r_out 500e-3
ri22 n141__r_out n143__r_out 500e-3
ri23 n155__r_out n153__r_out 500e-3
ri24 n154__r_out n156__r_out 500e-3
ri25 n168__r_out n158__r_out 500e-3
ri26 n159__r_out n169__r_out 500e-3
ri27 n174__r_out n171__r_out 500e-3
ri28 n172__r_out n175__r_out 500e-3
ri29 n194__r_out n184__r_out 500e-3
ri30 n185__r_out n195__r_out 500e-3
ri31 n200__r_out n197__r_out 500e-3
ri32 n198__r_out n201__r_out 500e-3
ri33 n220__r_out n218__r_out 500e-3
ri34 n219__r_out n221__r_out 500e-3
ri35 n226__r_out n223__r_out 500e-3
ri36 n224__r_out n227__r_out 500e-3
ri37 n239__r_out n236__r_out 500e-3
ri38 n237__r_out n240__r_out 500e-3
ri39 n252__r_out n249__r_out 500e-3
ri40 n250__r_out n253__r_out 500e-3
ri41 n265__r_out n262__r_out 500e-3
ri42 n263__r_out n266__r_out 500e-3
ri43 n285__r_out n283__r_out 500e-3
ri44 n284__r_out n286__r_out 500e-3
ri45 n291__r_out n288__r_out 500e-3
ri46 n289__r_out n292__r_out 500e-3
ri47 n304__r_out n301__r_out 500e-3
ri48 n302__r_out n305__r_out 500e-3
ri49 n317__r_out n314__r_out 500e-3
ri50 n315__r_out n318__r_out 500e-3
ri51 n330__r_out n327__r_out 500e-3
ri52 n328__r_out n331__r_out 500e-3
ri53 n350__r_out n348__r_out 500e-3
ri54 n349__r_out n351__r_out 500e-3
ri55 n363__r_out n353__r_out 500e-3
ri56 n354__r_out n364__r_out 500e-3
ri57 n369__r_out n366__r_out 500e-3
ri58 n367__r_out n370__r_out 500e-3
ri59 n389__r_out n379__r_out 500e-3
ri60 n380__r_out n390__r_out 500e-3
ri61 n402__r_out n392__r_out 500e-3
ri62 n393__r_out n403__r_out 500e-3
ri63 n415__r_out n413__r_out 500e-3
ri64 n414__r_out n416__r_out 500e-3
ri65 n428__r_out n426__r_out 500e-3
ri66 n427__r_out n429__r_out 500e-3
ri67 n436__r_out n433__r_out 500e-3
ri68 n434__r_out n437__r_out 500e-3
ri69 n456__r_out n454__r_out 500e-3
ri70 n455__r_out n457__r_out 500e-3
ri71 n472__r_out n470__r_out 500e-3
ri72 n471__r_out n473__r_out 500e-3
ri73 n485__r_out n475__r_out 500e-3
ri74 n476__r_out n486__r_out 500e-3
ri75 n491__r_out n488__r_out 500e-3
ri76 n489__r_out n492__r_out 500e-3
ri77 n5__x3 n4__x3 500e-3
ri78 n4__x2 n5__x2 500e-3
ri79 n5__x1 n4__x1 500e-3
ri80 n4__x0 n5__x0 500e-3
ri81 n12__reset n13__reset 1.1393
ri82 n14__reset n15__reset 1.9859
ri83 n8__i14__i17__net6 n9__i14__i17__net6 2.1908
ri84 n504__r_out n500__r_out 500e-3
ri85 n503__r_out n505__r_out 500e-3
ri86 n8__i14__i17__net1 n9__i14__i17__net1 1.2905
ri87 n4__i14__i17__net8 n5__i14__i17__net8 1.32
ri89 n12__i14__i17__net1 n13__i14__i17__net1 500e-3
ri90 n29__i14__net9 n21__i14__net9 1
ri91 n23__i14__net9 n30__i14__net9 1
ri92 n31__i14__net9 n25__i14__net9 1
ri93 n27__i14__net9 n32__i14__net9 1
ri94 n8__i14__i17__net7 n9__i14__i17__net7 1
ri95 n45__i14__net10 n37__i14__net10 1
ri96 n39__i14__net10 n46__i14__net10 1
ri97 n47__i14__net10 n41__i14__net10 1
ri98 n43__i14__net10 n48__i14__net10 1
ri99 n524__r_out n513__r_out 500e-3
ri100 n516__r_out n525__r_out 500e-3
ri101 n17__i14__net3 n9__i14__net3 500e-3
ri102 n12__i14__net3 n18__i14__net3 500e-3
ri103 n19__i14__net3 n13__i14__net3 500e-3
ri104 n16__i14__net3 n20__i14__net3 500e-3
ri105 n16__ck n19__ck 1
ri106 n537__r_out n535__r_out 500e-3
ri107 n536__r_out n538__r_out 500e-3
ri108 n25__reset n22__reset 1.0378
ri109 n550__r_out n548__r_out 500e-3
ri110 n549__r_out n551__r_out 500e-3
ri111 n563__r_out n561__r_out 500e-3
ri112 n562__r_out n564__r_out 500e-3
ri113 n2__vdd n7__vdd 83.33e-3
ri114 n8__vdd n3__vdd 83.33e-3
ri115 n6__vdd n9__vdd 83.33e-3
ri116 n9__i14__net4 n10__i14__net4 1
ri117 n11__i14__net4 n12__i14__net4 1
ri118 n13__i14__net4 n14__i14__net4 1
ri119 n15__i14__net4 n16__i14__net4 1
ri120 n576__r_out n574__r_out 500e-3
ri121 n575__r_out n577__r_out 500e-3
ri122 n13__i14__i17__net7 n14__i14__i17__net7 1.191
ri123 n587__r_out n588__r_out 1
ri124 n589__r_out n590__r_out 1
ri125 n21__i14__i17__net1 n22__i14__i17__net1 1.3265
ri130 n602__r_out n600__r_out 500e-3
ri131 n601__r_out n603__r_out 500e-3
ri132 n4__x_out_3 n5__x_out_3 790.3e-3
ri133 n5__x_out_2 n4__x_out_2 790.3e-3
ri134 n4__x_out_1 n5__x_out_1 790.3e-3
ri135 n5__x_out_0 n4__x_out_0 790.3e-3
ri136 n18__i14__i17__net8 n17__i14__i17__net8 766e-3
ri137 n23__i14__i17__net1 n24__i14__i17__net1 278.1e-3
ri138 n24__i14__i17__net1 n25__i14__i17__net1 894.8e-3
ri139 n4__y3 n5__y3 1.2817
ri140 n4__y2 n5__y2 1.2817
ri141 n4__y1 n5__y1 1.2817
ri142 n4__y0 n5__y0 1.2817
ri143 n15__i14__i17__net7 n16__i14__i17__net7 1.4311
ri144 n8__i14__i17__net11 n9__i14__i17__net11 1.3507
ri145 n615__r_out n613__r_out 500e-3
ri146 n614__r_out n616__r_out 500e-3
ri147 n10__i14__i17__net10 n8__i14__i17__net10 1.2581
ri148 n69__i14__net9 n61__i14__net9 1
ri149 n63__i14__net9 n70__i14__net9 1
ri150 n71__i14__net9 n65__i14__net9 1
ri151 n67__i14__net9 n72__i14__net9 1
ri152 n13__i14__i17__net9 n12__i14__i17__net9 1.3693
ri153 n628__r_out n626__r_out 500e-3
ri154 n627__r_out n629__r_out 500e-3
ri155 n89__i14__net10 n78__i14__net10 1
ri156 n79__i14__net10 n90__i14__net10 1
ri157 n91__i14__net10 n82__i14__net10 1
ri158 n83__i14__net10 n92__i14__net10 1
ri159 n46__reset n47__reset 1.685
ri160 n53__i14__net3 n49__i14__net3 500e-3
ri161 n50__i14__net3 n54__i14__net3 500e-3
ri162 n55__i14__net3 n51__i14__net3 500e-3
ri163 n52__i14__net3 n56__i14__net3 500e-3
ri164 n641__r_out n639__r_out 500e-3
ri165 n640__r_out n642__r_out 500e-3
ri166 n409__vss n401__vss 83.33e-3
ri167 n404__vss n410__vss 83.33e-3
ri168 n411__vss n405__vss 83.33e-3
ri169 n408__vss n412__vss 83.33e-3
ri170 n654__r_out n652__r_out 500e-3
ri171 n653__r_out n655__r_out 500e-3
ri173 n500__i18__net5 n498__i18__net5 127e-3
ri174 n498__i18__net5 n496__i18__net5 133.6e-3
ri175 n496__i18__net5 n494__i18__net5 137.4e-3
ri176 n494__i18__net5 n492__i18__net5 133.6e-3
ri177 n492__i18__net5 n490__i18__net5 129.8e-3
ri178 n490__i18__net5 n488__i18__net5 133.6e-3
ri179 n488__i18__net5 n486__i18__net5 133.6e-3
ri180 n486__i18__net5 n484__i18__net5 133.6e-3
ri181 n484__i18__net5 n482__i18__net5 133.6e-3
ri182 n482__i18__net5 n480__i18__net5 133.6e-3
ri183 n480__i18__net5 n478__i18__net5 133.6e-3
ri184 n478__i18__net5 n476__i18__net5 133.6e-3
ri185 n476__i18__net5 n474__i18__net5 137.4e-3
ri186 n474__i18__net5 n469__i18__net5 133.6e-3
ri187 n469__i18__net5 n466__i18__net5 129.8e-3
ri188 n466__i18__net5 n462__i18__net5 133.6e-3
ri189 n462__i18__net5 n457__i18__net5 133.6e-3
ri190 n457__i18__net5 n448__i18__net5 133.6e-3
ri191 n448__i18__net5 n447__i18__net5 133.6e-3
ri192 n447__i18__net5 n439__i18__net5 133.6e-3
ri193 n439__i18__net5 n433__i18__net5 133.6e-3
ri194 n433__i18__net5 n432__i18__net5 133.6e-3
ri195 n432__i18__net5 n427__i18__net5 137.4e-3
ri196 n427__i18__net5 n422__i18__net5 133.6e-3
ri197 n422__i18__net5 n417__i18__net5 129.8e-3
ri198 n417__i18__net5 n412__i18__net5 133.6e-3
ri199 n412__i18__net5 n404__i18__net5 133.6e-3
ri200 n404__i18__net5 n401__i18__net5 133.6e-3
ri201 n401__i18__net5 n394__i18__net5 133.6e-3
ri202 n394__i18__net5 n389__i18__net5 133.6e-3
ri203 n389__i18__net5 n384__i18__net5 133.6e-3
ri204 n384__i18__net5 n382__i18__net5 137.4e-3
ri205 n382__i18__net5 n374__i18__net5 133.6e-3
ri206 n374__i18__net5 n372__i18__net5 129.8e-3
ri207 n372__i18__net5 n364__i18__net5 133.6e-3
ri208 n364__i18__net5 n359__i18__net5 133.6e-3
ri209 n359__i18__net5 n354__i18__net5 133.6e-3
ri210 n354__i18__net5 n352__i18__net5 133.6e-3
ri211 n352__i18__net5 n344__i18__net5 133.6e-3
ri212 n344__i18__net5 n342__i18__net5 133.6e-3
ri213 n342__i18__net5 n334__i18__net5 133.6e-3
ri214 n334__i18__net5 n332__i18__net5 137.4e-3
ri215 n332__i18__net5 n324__i18__net5 133.6e-3
ri216 n324__i18__net5 n319__i18__net5 129.8e-3
ri217 n319__i18__net5 n317__i18__net5 133.6e-3
ri218 n317__i18__net5 n309__i18__net5 133.6e-3
ri219 n309__i18__net5 n307__i18__net5 133.6e-3
ri220 n307__i18__net5 n302__i18__net5 133.6e-3
ri221 n302__i18__net5 n297__i18__net5 133.6e-3
ri222 n297__i18__net5 n292__i18__net5 133.6e-3
ri223 n292__i18__net5 n287__i18__net5 133.6e-3
ri224 n287__i18__net5 n282__i18__net5 137.4e-3
ri225 n282__i18__net5 n274__i18__net5 133.6e-3
ri226 n274__i18__net5 n272__i18__net5 129.8e-3
ri227 n272__i18__net5 n264__i18__net5 133.6e-3
ri228 n264__i18__net5 n262__i18__net5 133.6e-3
ri229 n262__i18__net5 n257__i18__net5 133.6e-3
ri230 n257__i18__net5 n249__i18__net5 133.6e-3
ri231 n249__i18__net5 n244__i18__net5 133.6e-3
ri232 n244__i18__net5 n239__i18__net5 133.6e-3
ri233 n239__i18__net5 n234__i18__net5 137.4e-3
ri234 n234__i18__net5 n232__i18__net5 133.6e-3
ri235 n232__i18__net5 n227__i18__net5 129.8e-3
ri236 n227__i18__net5 n222__i18__net5 133.6e-3
ri237 n222__i18__net5 n217__i18__net5 133.6e-3
ri238 n217__i18__net5 n212__i18__net5 133.6e-3
ri239 n212__i18__net5 n207__i18__net5 133.6e-3
ri240 n207__i18__net5 n202__i18__net5 133.6e-3
ri241 n202__i18__net5 n197__i18__net5 133.6e-3
ri242 n197__i18__net5 n192__i18__net5 133.6e-3
ri243 n192__i18__net5 n184__i18__net5 137.4e-3
ri244 n184__i18__net5 n182__i18__net5 133.6e-3
ri245 n182__i18__net5 n177__i18__net5 129.8e-3
ri246 n177__i18__net5 n169__i18__net5 133.6e-3
ri247 n169__i18__net5 n167__i18__net5 133.6e-3
ri248 n167__i18__net5 n159__i18__net5 133.6e-3
ri249 n159__i18__net5 n157__i18__net5 133.6e-3
ri250 n157__i18__net5 n152__i18__net5 133.6e-3
ri251 n152__i18__net5 n147__i18__net5 133.6e-3
ri252 n147__i18__net5 n142__i18__net5 133.6e-3
ri253 n142__i18__net5 n134__i18__net5 137.4e-3
ri254 n134__i18__net5 n132__i18__net5 133.6e-3
ri255 n132__i18__net5 n127__i18__net5 129.8e-3
ri256 n127__i18__net5 n118__i18__net5 133.6e-3
ri257 n118__i18__net5 n114__i18__net5 133.6e-3
ri258 n114__i18__net5 n108__i18__net5 133.6e-3
ri259 n108__i18__net5 n107__i18__net5 133.6e-3
ri260 n107__i18__net5 n99__i18__net5 133.6e-3
ri261 n99__i18__net5 n94__i18__net5 133.6e-3
ri262 n94__i18__net5 n89__i18__net5 137.4e-3
ri263 n89__i18__net5 n84__i18__net5 133.6e-3
ri264 n84__i18__net5 n82__i18__net5 129.8e-3
ri265 n82__i18__net5 n77__i18__net5 133.6e-3
ri266 n77__i18__net5 n72__i18__net5 133.6e-3
ri267 n72__i18__net5 n67__i18__net5 133.6e-3
ri268 n67__i18__net5 n59__i18__net5 133.6e-3
ri269 n59__i18__net5 n57__i18__net5 133.6e-3
ri270 n57__i18__net5 n49__i18__net5 133.6e-3
ri271 n49__i18__net5 n47__i18__net5 133.6e-3
ri272 n58__i14__net4 n61__i14__net4 776e-3
ri273 n61__i14__net4 n62__i14__net4 491.2e-3
ri275 n62__i14__net4 n64__i14__net4 1.0072
ri277 n64__i14__net4 n66__i14__net4 388.1e-3
ri279 n66__i14__net4 n68__i14__net4 1.0072
ri280 n68__i14__net4 n69__i14__net4 500e-3
ri281 n29__i14__net11 n30__i14__net11 1.6089
ri282 n31__i14__net7 n32__i14__net7 1
ri283 n63__i14__net3 n64__i14__net3 952.8e-3
ri284 n64__i14__net3 n65__i14__net3 862.1e-3
ri285 n65__i14__net3 n66__i14__net3 533.2e-3
ri286 n66__i14__net3 n67__i14__net3 1.3621
ri287 n418__vddio n419__vddio 83.33e-3
ri288 n439__vss n433__vss 83.33e-3
ri289 n81__i14__net9 n82__i14__net9 1.8476
ri290 n82__i14__net9 n83__i14__net9 722.4e-3
ri291 n83__i14__net9 n84__i14__net9 678.3e-3
ri292 n84__i14__net9 n85__i14__net9 1.2224
ri293 n12__x_out_3 n13__x_out_3 1.2119
ri294 n12__x_out_2 n13__x_out_2 1.2119
ri295 n12__x_out_1 n13__x_out_1 1.2119
ri296 n10__x_out_0 n11__x_out_0 1.2119
ri301 n36__i14__net7 n35__i14__net7 500e-3
ri302 n33__i14__net11 n35__i14__net11 500e-3
ri303 n513__i18__net5 n503__i18__net5 500e-3
ri304 n504__i18__net5 n514__i18__net5 500e-3
ri309 n39__i14__net7 n38__i14__net7 500e-3
ri310 n37__i14__net11 n38__i14__net11 500e-3
ri311 n5__y_out_3 n6__y_out_3 1
ri312 n5__y_out_2 n6__y_out_2 1
ri313 n5__y_out_1 n6__y_out_1 1
ri314 n7__y_out_0 n8__y_out_0 1
ri315 n526__i18__net5 n524__i18__net5 500e-3
ri316 n525__i18__net5 n527__i18__net5 500e-3
ri317 n106__i14__net10 n109__i14__net10 679.1e-3
ri318 n109__i14__net10 n110__i14__net10 426.8e-3
ri319 n110__i14__net10 n111__i14__net10 985.7e-3
ri320 n111__i14__net10 n112__i14__net10 926.8e-3
ri321 n14__x_out_2 n15__x_out_2 1
ri322 n12__y_out_0 n13__y_out_0 1
ri323 n12__x_out_0 n13__x_out_0 1
ri324 n10__y_out_2 n11__y_out_2 1
ri325 n539__i18__net5 n537__i18__net5 500e-3
ri326 n538__i18__net5 n540__i18__net5 500e-3
ri327 n19__x_out_2 n20__x_out_2 1.652
ri328 n15__y_out_2 n16__y_out_2 1.6762
ri329 n552__i18__net5 n550__i18__net5 500e-3
ri330 n551__i18__net5 n553__i18__net5 500e-3
ri331 n14__ck_b n12__ck_b 628.8e-3
ri332 n12__ck_b n15__ck_b 818e-3
ri333 n8__ck_buff n9__ck_buff 1.3446
ri334 n3__reset_b n4__reset_b 1.3343
ri335 n5__reset_b n6__reset_b 1
ri336 n558__i18__net5 n555__i18__net5 500e-3
ri337 n556__i18__net5 n559__i18__net5 500e-3
ri338 n19__i13__a2 n20__i13__a2 1.2672
ri339 n19__i13__a0 n20__i13__a0 1.2672
ri340 n7__reset_buff n6__reset_buff 500e-3
ri341 n14__x_out_3 n15__x_out_3 1.8603
ri343 n14__x_out_1 n15__x_out_1 1
ri344 n576__i18__net5 n578__i18__net5 500e-3
ri345 n579__i18__net5 n577__i18__net5 500e-3
ri346 n8__reset_buff n9__reset_buff 1.4607
ri347 n10__y_out_1 n11__y_out_1 1
ri348 n10__y_out_3 n11__y_out_3 2.0514
ri349 n11__y_out_3 n12__y_out_3 500e-3
ri350 n30__ck n32__ck 1.185
ri351 n15__y_out_1 n16__y_out_1 2.1886
ri352 n20__x_out_1 n21__x_out_1 2.0356
ri353 n591__i18__net5 n589__i18__net5 500e-3
ri354 n590__i18__net5 n592__i18__net5 500e-3
ri355 n597__i18__net5 n594__i18__net5 500e-3
ri356 n595__i18__net5 n598__i18__net5 500e-3
ri357 n21__i13__a2 n22__i13__a2 1.0883
ri358 n18__i13__a3 n17__i13__a3 573.7e-3
ri359 n17__i13__a1 n18__i13__a1 573.7e-3
ri360 n21__i13__a0 n22__i13__a0 1.0883
ri361 n507__vss n504__vss 83.33e-3
ri362 n505__vss n508__vss 83.33e-3
ri363 n35__ck n36__ck 250e-3
ri364 n617__i18__net5 n615__i18__net5 500e-3
ri365 n616__i18__net5 n618__i18__net5 500e-3
ri366 n61__reset n62__reset 250e-3
ri367 n628__i18__net5 n630__i18__net5 500e-3
ri368 n631__i18__net5 n629__i18__net5 500e-3
ri369 n64__reset n65__reset 250e-3
ri370 n22__ck_buff n23__ck_buff 1.1753
ri371 n632__i18__net5 n633__i18__net5 1
ri372 n634__i18__net5 n635__i18__net5 1
ri373 r0_buff n2__r0_buff 2.3911
ri374 n654__i18__net5 n656__i18__net5 500e-3
ri375 n657__i18__net5 n655__i18__net5 500e-3
ri376 n17__ck4 n9__ck4 3.1516
ri377 n9__ck4 n5__ck4 656.2e-3
ri378 r1_buff n2__r1_buff 1.6061
ri380 n16__reset_buff n19__reset_buff 653e-3
ri381 r2_buff n2__r2_buff 1.4196
ri382 n17__i13__net12 n18__i13__net12 1.544
ri383 n15__i13__net1 n16__i13__net1 2.0685
ri384 n669__i18__net5 n667__i18__net5 500e-3
ri385 n668__i18__net5 n670__i18__net5 500e-3
ri386 n13__i13__net11 n14__i13__net11 745.7e-3
ri387 n19__i13__net2 n20__i13__net2 673.2e-3
ri388 n3__net3 n2__net3 934.5e-3
ri389 net4 n3__net4 513.2e-3
ri390 n531__vss n526__vss 394e-3
ri391 n675__i18__net5 n671__i18__net5 500e-3
ri392 n674__i18__net5 n676__i18__net5 500e-3
ri393 n6__r0_buff n7__r0_buff 897.8e-3
ri394 n6__r1_buff n7__r1_buff 784.9e-3
ri395 n6__r2_buff n7__r2_buff 697.9e-3
ri396 n25__vdd n24__vdd 83.33e-3
ri397 n6__net4 n7__net4 1.315
ri398 n693__i18__net5 n695__i18__net5 500e-3
ri399 n696__i18__net5 n694__i18__net5 500e-3
ri400 n31__ck_b n32__ck_b 873.6e-3
ri401 n32__ck_b n33__ck_b 699.3e-3
ri402 n33__ck_b n34__ck_b 1.2346
ri404 n150__i18__net4 n148__i18__net4 127e-3
ri405 n148__i18__net4 n146__i18__net4 133.6e-3
ri406 n146__i18__net4 n144__i18__net4 137.4e-3
ri407 n144__i18__net4 n142__i18__net4 133.6e-3
ri408 n142__i18__net4 n140__i18__net4 129.8e-3
ri409 n140__i18__net4 n138__i18__net4 133.6e-3
ri410 n138__i18__net4 n136__i18__net4 133.6e-3
ri411 n136__i18__net4 n134__i18__net4 133.6e-3
ri412 n134__i18__net4 n132__i18__net4 133.6e-3
ri413 n132__i18__net4 n130__i18__net4 133.6e-3
ri414 n130__i18__net4 n128__i18__net4 133.6e-3
ri415 n128__i18__net4 n126__i18__net4 133.6e-3
ri416 n126__i18__net4 n124__i18__net4 137.4e-3
ri417 n124__i18__net4 n118__i18__net4 133.6e-3
ri418 n118__i18__net4 n117__i18__net4 129.8e-3
ri419 n117__i18__net4 n109__i18__net4 133.6e-3
ri420 n109__i18__net4 n107__i18__net4 133.6e-3
ri421 n107__i18__net4 n99__i18__net4 133.6e-3
ri422 n99__i18__net4 n93__i18__net4 133.6e-3
ri423 n93__i18__net4 n92__i18__net4 133.6e-3
ri424 n92__i18__net4 n87__i18__net4 133.6e-3
ri425 n87__i18__net4 n79__i18__net4 133.6e-3
ri426 n79__i18__net4 n77__i18__net4 137.4e-3
ri427 n77__i18__net4 n72__i18__net4 133.6e-3
ri428 n72__i18__net4 n67__i18__net4 129.8e-3
ri429 n67__i18__net4 n62__i18__net4 133.6e-3
ri430 n62__i18__net4 n57__i18__net4 133.6e-3
ri431 n57__i18__net4 n52__i18__net4 133.6e-3
ri432 n52__i18__net4 n44__i18__net4 133.6e-3
ri433 n26__reset_buff n27__reset_buff 1.0597
ri434 n27__reset_buff n28__reset_buff 65.86e-3
ri435 n28__reset_buff n29__reset_buff 1.3314
ri436 n34__ck_buff n35__ck_buff 947.7e-3
ri437 n34__ck_buff n36__ck_buff 1.0268
ri438 n36__ck_buff n37__ck_buff 850.9e-3
ri439 n21__reset_b n22__reset_b 939.6e-3
ri440 n22__reset_b n23__reset_b 397.3e-3
ri441 n23__reset_b n24__reset_b 1.5317
ri442 n161__i18__net4 n159__i18__net4 500e-3
ri443 n160__i18__net4 n162__i18__net4 500e-3
ri444 n21__i13__net18 n19__i13__net18 679e-3
ri445 n13__i13__net7 n15__i13__net7 1.3877
ri446 n10__i13__net17 n11__i13__net17 964.9e-3
ri447 n172__i18__net4 n170__i18__net4 500e-3
ri448 n171__i18__net4 n173__i18__net4 500e-3
ri449 n174__i18__net4 n175__i18__net4 1
ri450 n176__i18__net4 n177__i18__net4 1
ri451 n11__i13__net23 n10__i13__net23 1.5439
ri452 n194__i18__net4 n192__i18__net4 500e-3
ri453 n193__i18__net4 n195__i18__net4 500e-3
ri454 n205__i18__net4 n203__i18__net4 500e-3
ri455 n204__i18__net4 n206__i18__net4 500e-3
ri456 n50__i18__net3 n48__i18__net3 133.6e-3
ri457 n48__i18__net3 n47__i18__net3 137.4e-3
ri458 n47__i18__net3 n44__i18__net3 133.6e-3
ri459 n44__i18__net3 n42__i18__net3 129.8e-3
ri460 n42__i18__net3 n40__i18__net3 133.6e-3
ri461 n40__i18__net3 n38__i18__net3 133.6e-3
ri462 n38__i18__net3 n37__i18__net3 133.6e-3
ri463 n37__i18__net3 n34__i18__net3 133.6e-3
ri464 n34__i18__net3 n32__i18__net3 133.6e-3
ri465 n14__serial_out_b_high n16__serial_out_b_high 1
ri466 n25__serial_out n29__serial_out 500e-3
ri469 n17__net4 n16__net4 500e-3
ri470 n14__net3 n15__net3 500e-3
ri472 n30__serial_out n26__serial_out 2.4328
ri473 n15__r1 n8__r1 3.163
ri474 n15__r0 n9__r0 5.82
ri475 n10__r2 n4__r2 4.56
ri476 n419__vdd n421__vdd 83.33e-3
ri477 n422__vdd n420__vdd 83.33e-3
ri478 n31__serial_out n32__serial_out 2.9745
ri479 n15__serial_out_b_high n17__serial_out_b_high 500e-3
ri480 n976__vddio n969__vddio 83.33e-3
ri481 n970__vddio n977__vddio 83.33e-3
ri482 n978__vddio n975__vddio 83.33e-3
ri483 n16__r0_buff n15__r0_buff 500e-3
ri484 n16__r2_buff n17__r2_buff 500e-3
ri485 n16__r1_buff n15__r1_buff 500e-3
ri486 n1304__vss n1309__vss 83.33e-3
ri488 n1308__vss n1303__vss 355.9e-3
ri489 n1303__vss n614__vss 1.4469
ri490 n614__vss n438__vss 2.1001
ri492 n438__vss n424__vss 128.3e-3
ri493 n424__vss n400__vss 120e-3
ri494 n400__vss n391__vss 124.6e-3
ri495 n391__vss n384__vss 133e-3
ri496 n384__vss n376__vss 124.6e-3
ri497 n376__vss n368__vss 124.6e-3
ri498 n368__vss n360__vss 124.6e-3
ri499 n360__vss n351__vss 120e-3
ri500 n351__vss n344__vss 124.6e-3
ri501 n344__vss n336__vss 133e-3
ri502 n336__vss n328__vss 124.6e-3
ri503 n328__vss n320__vss 120e-3
ri504 n320__vss n312__vss 124.6e-3
ri505 n312__vss n304__vss 125.5e-3
ri506 n304__vss n296__vss 124.6e-3
ri507 n296__vss n288__vss 120e-3
ri508 n288__vss n280__vss 124.6e-3
ri509 n280__vss n272__vss 133e-3
ri510 n272__vss n264__vss 124.6e-3
ri511 n264__vss n256__vss 120e-3
ri512 n256__vss n248__vss 125.5e-3
ri513 n248__vss n240__vss 124.6e-3
ri514 n240__vss n232__vss 120e-3
ri515 n232__vss n224__vss 124.6e-3
ri516 n224__vss n216__vss 133e-3
ri517 n216__vss n208__vss 124.6e-3
ri518 n208__vss n200__vss 120e-3
ri519 n200__vss n192__vss 124.6e-3
ri520 n192__vss n184__vss 125.5e-3
ri521 n184__vss n176__vss 124.6e-3
ri522 n176__vss n168__vss 120e-3
ri523 n168__vss n160__vss 124.6e-3
ri524 n160__vss n152__vss 133e-3
ri525 n152__vss n144__vss 124.6e-3
ri526 n144__vss n136__vss 120e-3
ri527 n136__vss n128__vss 121.8e-3
ri528 n128__vss n120__vss 124.6e-3
ri529 n120__vss n112__vss 120e-3
ri530 n112__vss n104__vss 124.6e-3
ri531 n104__vss n96__vss 133e-3
ri532 n96__vss n88__vss 124.6e-3
ri533 n88__vss n80__vss 120e-3
ri534 n80__vss n72__vss 124.6e-3
ri535 n72__vss n64__vss 125.5e-3
ri536 n64__vss n56__vss 124.6e-3
ri537 n56__vss n48__vss 120e-3
ri538 n48__vss n40__vss 124.6e-3
ri539 n40__vss n32__vss 133e-3
ri540 n32__vss n24__vss 124.6e-3
ri541 n24__vss n16__vss 120e-3
ri542 n16__vss n8__vss 124.6e-3
ri544 n971__vddio n968__vddio 169.1e-3
ri545 n968__vddio n633__vddio 1.4469
ri546 n633__vddio n530__vddio 124.6e-3
ri547 n530__vddio n524__vddio 133e-3
ri548 n524__vddio n518__vddio 124.6e-3
ri549 n518__vddio n512__vddio 124.6e-3
ri550 n512__vddio n505__vddio 124.6e-3
ri551 n505__vddio n499__vddio 120e-3
ri552 n499__vddio n494__vddio 124.6e-3
ri553 n494__vddio n488__vddio 133e-3
ri554 n488__vddio n482__vddio 124.6e-3
ri555 n482__vddio n476__vddio 120e-3
ri556 n476__vddio n470__vddio 111.6e-3
ri557 n470__vddio n464__vddio 124.6e-3
ri558 n464__vddio n457__vddio 133e-3
ri559 n457__vddio n451__vddio 124.6e-3
ri560 n451__vddio n430__vddio 120e-3
ri561 n430__vddio n413__vddio 152.7e-3
ri563 n413__vddio n401__vddio 124.8e-3
ri564 n401__vddio n393__vddio 120e-3
ri565 n393__vddio n386__vddio 124.6e-3
ri566 n386__vddio n377__vddio 133e-3
ri567 n377__vddio n369__vddio 124.6e-3
ri568 n369__vddio n361__vddio 124.6e-3
ri569 n361__vddio n353__vddio 124.6e-3
ri570 n353__vddio n346__vddio 120e-3
ri571 n346__vddio n337__vddio 124.6e-3
ri572 n337__vddio n329__vddio 133e-3
ri573 n329__vddio n321__vddio 124.6e-3
ri574 n321__vddio n313__vddio 120e-3
ri575 n313__vddio n305__vddio 124.6e-3
ri576 n305__vddio n297__vddio 125.5e-3
ri577 n297__vddio n289__vddio 124.6e-3
ri578 n289__vddio n281__vddio 120e-3
ri579 n281__vddio n273__vddio 124.6e-3
ri580 n273__vddio n265__vddio 133e-3
ri581 n265__vddio n257__vddio 124.6e-3
ri582 n257__vddio n249__vddio 120e-3
ri583 n249__vddio n241__vddio 125.5e-3
ri584 n241__vddio n233__vddio 124.6e-3
ri585 n233__vddio n225__vddio 120e-3
ri586 n225__vddio n217__vddio 124.6e-3
ri587 n217__vddio n209__vddio 133e-3
ri588 n209__vddio n201__vddio 124.6e-3
ri589 n201__vddio n193__vddio 120e-3
ri590 n193__vddio n185__vddio 124.6e-3
ri591 n185__vddio n177__vddio 125.5e-3
ri592 n177__vddio n169__vddio 124.6e-3
ri593 n169__vddio n161__vddio 120e-3
ri594 n161__vddio n153__vddio 124.6e-3
ri595 n153__vddio n145__vddio 133e-3
ri596 n145__vddio n137__vddio 124.6e-3
ri597 n137__vddio n129__vddio 120e-3
ri598 n129__vddio n121__vddio 121.8e-3
ri599 n121__vddio n113__vddio 124.6e-3
ri600 n113__vddio n105__vddio 120e-3
ri601 n105__vddio n97__vddio 124.6e-3
ri602 n97__vddio n89__vddio 133e-3
ri603 n89__vddio n81__vddio 124.6e-3
ri604 n81__vddio n73__vddio 120e-3
ri605 n73__vddio n65__vddio 124.6e-3
ri606 n65__vddio n57__vddio 125.5e-3
ri607 n57__vddio n49__vddio 124.6e-3
ri608 n49__vddio n41__vddio 120e-3
ri609 n41__vddio n33__vddio 124.6e-3
ri610 n33__vddio n25__vddio 133e-3
ri611 n25__vddio n17__vddio 124.6e-3
ri612 n17__vddio n9__vddio 120e-3
ri613 n9__vddio n1__vddio 124.6e-3
ri615 n972__vddio n967__vddio 493.4e-3
ri616 n967__vddio n634__vddio 1.1226
ri617 n634__vddio n531__vddio 124.6e-3
ri618 n531__vddio n525__vddio 133e-3
ri619 n525__vddio n519__vddio 124.6e-3
ri620 n519__vddio n513__vddio 124.6e-3
ri621 n513__vddio n508__vddio 124.6e-3
ri622 n508__vddio n502__vddio 120e-3
ri623 n502__vddio n495__vddio 124.6e-3
ri624 n495__vddio n489__vddio 133e-3
ri625 n489__vddio n483__vddio 124.6e-3
ri626 n483__vddio n477__vddio 120e-3
ri627 n477__vddio n471__vddio 111.6e-3
ri628 n471__vddio n465__vddio 124.6e-3
ri629 n465__vddio n460__vddio 133e-3
ri630 n460__vddio n454__vddio 124.6e-3
ri631 n454__vddio n431__vddio 120e-3
ri632 n431__vddio n414__vddio 153.4e-3
ri634 n414__vddio n404__vddio 125.5e-3
ri635 n404__vddio n396__vddio 120e-3
ri636 n396__vddio n387__vddio 124.6e-3
ri637 n387__vddio n380__vddio 133e-3
ri638 n380__vddio n372__vddio 124.6e-3
ri639 n372__vddio n364__vddio 124.6e-3
ri640 n364__vddio n356__vddio 124.6e-3
ri641 n356__vddio n347__vddio 120e-3
ri642 n347__vddio n340__vddio 124.6e-3
ri643 n340__vddio n332__vddio 133e-3
ri644 n332__vddio n324__vddio 124.6e-3
ri645 n324__vddio n316__vddio 120e-3
ri646 n316__vddio n308__vddio 124.6e-3
ri647 n308__vddio n300__vddio 125.5e-3
ri648 n300__vddio n292__vddio 124.6e-3
ri649 n292__vddio n284__vddio 120e-3
ri650 n284__vddio n276__vddio 124.6e-3
ri651 n276__vddio n268__vddio 133e-3
ri652 n268__vddio n260__vddio 124.6e-3
ri653 n260__vddio n252__vddio 120e-3
ri654 n252__vddio n244__vddio 125.5e-3
ri655 n244__vddio n236__vddio 124.6e-3
ri656 n236__vddio n228__vddio 120e-3
ri657 n228__vddio n220__vddio 124.6e-3
ri658 n220__vddio n212__vddio 133e-3
ri659 n212__vddio n204__vddio 124.6e-3
ri660 n204__vddio n196__vddio 120e-3
ri661 n196__vddio n188__vddio 124.6e-3
ri662 n188__vddio n180__vddio 125.5e-3
ri663 n180__vddio n172__vddio 124.6e-3
ri664 n172__vddio n164__vddio 120e-3
ri665 n164__vddio n156__vddio 124.6e-3
ri666 n156__vddio n148__vddio 133e-3
ri667 n148__vddio n140__vddio 124.6e-3
ri668 n140__vddio n132__vddio 120e-3
ri669 n132__vddio n124__vddio 121.8e-3
ri670 n124__vddio n116__vddio 124.6e-3
ri671 n116__vddio n108__vddio 120e-3
ri672 n108__vddio n100__vddio 124.6e-3
ri673 n100__vddio n92__vddio 133e-3
ri674 n92__vddio n84__vddio 124.6e-3
ri675 n84__vddio n76__vddio 120e-3
ri676 n76__vddio n68__vddio 124.6e-3
ri677 n68__vddio n60__vddio 125.5e-3
ri678 n60__vddio n52__vddio 124.6e-3
ri679 n52__vddio n44__vddio 120e-3
ri680 n44__vddio n36__vddio 124.6e-3
ri681 n36__vddio n28__vddio 133e-3
ri682 n28__vddio n20__vddio 124.6e-3
ri683 n20__vddio n12__vddio 120e-3
ri684 n12__vddio n4__vddio 124.6e-3
ri686 n973__vddio n982__vddio 829.8e-3
ri687 n982__vddio n983__vddio 338.2e-3
ri688 n983__vddio n635__vddio 447.9e-3
ri689 n635__vddio n534__vddio 124.6e-3
ri690 n534__vddio n528__vddio 133e-3
ri691 n528__vddio n522__vddio 124.6e-3
ri692 n522__vddio n516__vddio 124.6e-3
ri693 n516__vddio n509__vddio 124.6e-3
ri694 n509__vddio n503__vddio 120e-3
ri695 n503__vddio n498__vddio 124.6e-3
ri696 n498__vddio n492__vddio 133e-3
ri697 n492__vddio n486__vddio 124.6e-3
ri698 n486__vddio n480__vddio 120e-3
ri699 n480__vddio n474__vddio 111.6e-3
ri700 n474__vddio n468__vddio 124.6e-3
ri701 n468__vddio n461__vddio 133e-3
ri702 n461__vddio n455__vddio 124.6e-3
ri703 n455__vddio n434__vddio 120e-3
ri704 n434__vddio n415__vddio 153.4e-3
ri706 n415__vddio n405__vddio 125.5e-3
ri707 n405__vddio n397__vddio 120e-3
ri708 n397__vddio n390__vddio 124.6e-3
ri709 n390__vddio n381__vddio 133e-3
ri710 n381__vddio n373__vddio 124.6e-3
ri711 n373__vddio n365__vddio 124.6e-3
ri712 n365__vddio n357__vddio 124.6e-3
ri713 n357__vddio n350__vddio 120e-3
ri714 n350__vddio n341__vddio 124.6e-3
ri715 n341__vddio n333__vddio 133e-3
ri716 n333__vddio n325__vddio 124.6e-3
ri717 n325__vddio n317__vddio 120e-3
ri718 n317__vddio n309__vddio 124.6e-3
ri719 n309__vddio n301__vddio 125.5e-3
ri720 n301__vddio n293__vddio 124.6e-3
ri721 n293__vddio n285__vddio 120e-3
ri722 n285__vddio n277__vddio 124.6e-3
ri723 n277__vddio n269__vddio 133e-3
ri724 n269__vddio n261__vddio 124.6e-3
ri725 n261__vddio n253__vddio 120e-3
ri726 n253__vddio n245__vddio 125.5e-3
ri727 n245__vddio n237__vddio 124.6e-3
ri728 n237__vddio n229__vddio 120e-3
ri729 n229__vddio n221__vddio 124.6e-3
ri730 n221__vddio n213__vddio 133e-3
ri731 n213__vddio n205__vddio 124.6e-3
ri732 n205__vddio n197__vddio 120e-3
ri733 n197__vddio n189__vddio 124.6e-3
ri734 n189__vddio n181__vddio 125.5e-3
ri735 n181__vddio n173__vddio 124.6e-3
ri736 n173__vddio n165__vddio 120e-3
ri737 n165__vddio n157__vddio 124.6e-3
ri738 n157__vddio n149__vddio 133e-3
ri739 n149__vddio n141__vddio 124.6e-3
ri740 n141__vddio n133__vddio 120e-3
ri741 n133__vddio n125__vddio 121.8e-3
ri742 n125__vddio n117__vddio 124.6e-3
ri743 n117__vddio n109__vddio 120e-3
ri744 n109__vddio n101__vddio 124.6e-3
ri745 n101__vddio n93__vddio 133e-3
ri746 n93__vddio n85__vddio 124.6e-3
ri747 n85__vddio n77__vddio 120e-3
ri748 n77__vddio n69__vddio 124.6e-3
ri749 n69__vddio n61__vddio 125.5e-3
ri750 n61__vddio n53__vddio 124.6e-3
ri751 n53__vddio n45__vddio 120e-3
ri752 n45__vddio n37__vddio 124.6e-3
ri753 n37__vddio n29__vddio 133e-3
ri754 n29__vddio n21__vddio 124.6e-3
ri755 n21__vddio n13__vddio 120e-3
ri756 n13__vddio n5__vddio 124.6e-3
ri757 n964__vddio n982__vddio 83.33e-3
ri758 n966__vddio n983__vddio 25e-3
ri760 n1305__vss n1312__vss 2.0034
ri761 n1312__vss n1313__vss 468.3e-3
ri762 n1313__vss n1314__vss 520.4e-3
ri763 n1314__vss n613__vss 520.4e-3
ri764 n613__vss n435__vss 395.9e-3
ri766 n435__vss n417__vss 128.3e-3
ri767 n417__vss n393__vss 120e-3
ri768 n393__vss n386__vss 124.6e-3
ri769 n386__vss n377__vss 133e-3
ri770 n377__vss n369__vss 124.6e-3
ri771 n369__vss n361__vss 124.6e-3
ri772 n361__vss n353__vss 124.6e-3
ri773 n353__vss n346__vss 120e-3
ri774 n346__vss n337__vss 124.6e-3
ri775 n337__vss n329__vss 133e-3
ri776 n329__vss n321__vss 124.6e-3
ri777 n321__vss n313__vss 120e-3
ri778 n313__vss n305__vss 124.6e-3
ri779 n305__vss n297__vss 125.5e-3
ri780 n297__vss n289__vss 124.6e-3
ri781 n289__vss n281__vss 120e-3
ri782 n281__vss n273__vss 124.6e-3
ri783 n273__vss n265__vss 133e-3
ri784 n265__vss n257__vss 124.6e-3
ri785 n257__vss n249__vss 120e-3
ri786 n249__vss n241__vss 125.5e-3
ri787 n241__vss n233__vss 124.6e-3
ri788 n233__vss n225__vss 120e-3
ri789 n225__vss n217__vss 124.6e-3
ri790 n217__vss n209__vss 133e-3
ri791 n209__vss n201__vss 124.6e-3
ri792 n201__vss n193__vss 120e-3
ri793 n193__vss n185__vss 124.6e-3
ri794 n185__vss n177__vss 125.5e-3
ri795 n177__vss n169__vss 124.6e-3
ri796 n169__vss n161__vss 120e-3
ri797 n161__vss n153__vss 124.6e-3
ri798 n153__vss n145__vss 133e-3
ri799 n145__vss n137__vss 124.6e-3
ri800 n137__vss n129__vss 120e-3
ri801 n129__vss n121__vss 121.8e-3
ri802 n121__vss n113__vss 124.6e-3
ri803 n113__vss n105__vss 120e-3
ri804 n105__vss n97__vss 124.6e-3
ri805 n97__vss n89__vss 133e-3
ri806 n89__vss n81__vss 124.6e-3
ri807 n81__vss n73__vss 120e-3
ri808 n73__vss n65__vss 124.6e-3
ri809 n65__vss n57__vss 125.5e-3
ri810 n57__vss n49__vss 124.6e-3
ri811 n49__vss n41__vss 120e-3
ri812 n41__vss n33__vss 124.6e-3
ri813 n33__vss n25__vss 133e-3
ri814 n25__vss n17__vss 124.6e-3
ri815 n17__vss n9__vss 120e-3
ri816 n9__vss n1__vss 124.6e-3
ri817 n606__vss n1312__vss 31.25e-3
ri818 n608__vss n1313__vss 25e-3
ri819 n610__vss n1314__vss 25e-3
ri821 n1306__vss n1316__vss 1.0166
ri822 n1316__vss n1301__vss 338.2e-3
ri823 n1301__vss n436__vss 2.5535
ri825 n436__vss n420__vss 128.3e-3
ri826 n420__vss n396__vss 120e-3
ri827 n396__vss n387__vss 124.6e-3
ri828 n387__vss n380__vss 133e-3
ri829 n380__vss n372__vss 124.6e-3
ri830 n372__vss n364__vss 124.6e-3
ri831 n364__vss n356__vss 124.6e-3
ri832 n356__vss n347__vss 120e-3
ri833 n347__vss n340__vss 124.6e-3
ri834 n340__vss n332__vss 133e-3
ri835 n332__vss n324__vss 124.6e-3
ri836 n324__vss n316__vss 120e-3
ri837 n316__vss n308__vss 124.6e-3
ri838 n308__vss n300__vss 125.5e-3
ri839 n300__vss n292__vss 124.6e-3
ri840 n292__vss n284__vss 120e-3
ri841 n284__vss n276__vss 124.6e-3
ri842 n276__vss n268__vss 133e-3
ri843 n268__vss n260__vss 124.6e-3
ri844 n260__vss n252__vss 120e-3
ri845 n252__vss n244__vss 125.5e-3
ri846 n244__vss n236__vss 124.6e-3
ri847 n236__vss n228__vss 120e-3
ri848 n228__vss n220__vss 124.6e-3
ri849 n220__vss n212__vss 133e-3
ri850 n212__vss n204__vss 124.6e-3
ri851 n204__vss n196__vss 120e-3
ri852 n196__vss n188__vss 124.6e-3
ri853 n188__vss n180__vss 125.5e-3
ri854 n180__vss n172__vss 124.6e-3
ri855 n172__vss n164__vss 120e-3
ri856 n164__vss n156__vss 124.6e-3
ri857 n156__vss n148__vss 133e-3
ri858 n148__vss n140__vss 124.6e-3
ri859 n140__vss n132__vss 120e-3
ri860 n132__vss n124__vss 121.8e-3
ri861 n124__vss n116__vss 124.6e-3
ri862 n116__vss n108__vss 120e-3
ri863 n108__vss n100__vss 124.6e-3
ri864 n100__vss n92__vss 133e-3
ri865 n92__vss n84__vss 124.6e-3
ri866 n84__vss n76__vss 120e-3
ri867 n76__vss n68__vss 124.6e-3
ri868 n68__vss n60__vss 125.5e-3
ri869 n60__vss n52__vss 124.6e-3
ri870 n52__vss n44__vss 120e-3
ri871 n44__vss n36__vss 124.6e-3
ri872 n36__vss n28__vss 133e-3
ri873 n28__vss n20__vss 124.6e-3
ri874 n20__vss n12__vss 120e-3
ri875 n12__vss n4__vss 124.6e-3
ri876 n1298__vss n1316__vss 83.33e-3
ri878 n1307__vss n1302__vss 680.2e-3
ri879 n1302__vss n437__vss 3.2281
ri881 n437__vss n421__vss 128.3e-3
ri882 n421__vss n397__vss 120e-3
ri883 n397__vss n390__vss 124.6e-3
ri884 n390__vss n381__vss 133e-3
ri885 n381__vss n373__vss 124.6e-3
ri886 n373__vss n365__vss 124.6e-3
ri887 n365__vss n357__vss 124.6e-3
ri888 n357__vss n350__vss 120e-3
ri889 n350__vss n341__vss 124.6e-3
ri890 n341__vss n333__vss 133e-3
ri891 n333__vss n325__vss 124.6e-3
ri892 n325__vss n317__vss 120e-3
ri893 n317__vss n309__vss 124.6e-3
ri894 n309__vss n301__vss 125.5e-3
ri895 n301__vss n293__vss 124.6e-3
ri896 n293__vss n285__vss 120e-3
ri897 n285__vss n277__vss 124.6e-3
ri898 n277__vss n269__vss 133e-3
ri899 n269__vss n261__vss 124.6e-3
ri900 n261__vss n253__vss 120e-3
ri901 n253__vss n245__vss 125.5e-3
ri902 n245__vss n237__vss 124.6e-3
ri903 n237__vss n229__vss 120e-3
ri904 n229__vss n221__vss 124.6e-3
ri905 n221__vss n213__vss 133e-3
ri906 n213__vss n205__vss 124.6e-3
ri907 n205__vss n197__vss 120e-3
ri908 n197__vss n189__vss 124.6e-3
ri909 n189__vss n181__vss 125.5e-3
ri910 n181__vss n173__vss 124.6e-3
ri911 n173__vss n165__vss 120e-3
ri912 n165__vss n157__vss 124.6e-3
ri913 n157__vss n149__vss 133e-3
ri914 n149__vss n141__vss 124.6e-3
ri915 n141__vss n133__vss 120e-3
ri916 n133__vss n125__vss 121.8e-3
ri917 n125__vss n117__vss 124.6e-3
ri918 n117__vss n109__vss 120e-3
ri919 n109__vss n101__vss 124.6e-3
ri920 n101__vss n93__vss 133e-3
ri921 n93__vss n85__vss 124.6e-3
ri922 n85__vss n77__vss 120e-3
ri923 n77__vss n69__vss 124.6e-3
ri924 n69__vss n61__vss 125.5e-3
ri925 n61__vss n53__vss 124.6e-3
ri926 n53__vss n45__vss 120e-3
ri927 n45__vss n37__vss 124.6e-3
ri928 n37__vss n29__vss 133e-3
ri929 n29__vss n21__vss 124.6e-3
ri930 n21__vss n13__vss 120e-3
ri931 n13__vss n5__vss 124.6e-3
ri933 n974__vddio n985__vddio 1.8166
ri934 n985__vddio n986__vddio 468.3e-3
ri935 n986__vddio n987__vddio 520.4e-3
ri936 n987__vddio n988__vddio 520.4e-3
ri937 n988__vddio n416__vddio 398.6e-3
ri939 n416__vddio n408__vddio 125.5e-3
ri940 n408__vddio n400__vddio 120e-3
ri941 n400__vddio n391__vddio 124.6e-3
ri942 n391__vddio n384__vddio 133e-3
ri943 n384__vddio n376__vddio 124.6e-3
ri944 n376__vddio n368__vddio 124.6e-3
ri945 n368__vddio n360__vddio 124.6e-3
ri946 n360__vddio n351__vddio 120e-3
ri947 n351__vddio n344__vddio 124.6e-3
ri948 n344__vddio n336__vddio 133e-3
ri949 n336__vddio n328__vddio 124.6e-3
ri950 n328__vddio n320__vddio 120e-3
ri951 n320__vddio n312__vddio 124.6e-3
ri952 n312__vddio n304__vddio 125.5e-3
ri953 n304__vddio n296__vddio 124.6e-3
ri954 n296__vddio n288__vddio 120e-3
ri955 n288__vddio n280__vddio 124.6e-3
ri956 n280__vddio n272__vddio 133e-3
ri957 n272__vddio n264__vddio 124.6e-3
ri958 n264__vddio n256__vddio 120e-3
ri959 n256__vddio n248__vddio 125.5e-3
ri960 n248__vddio n240__vddio 124.6e-3
ri961 n240__vddio n232__vddio 120e-3
ri962 n232__vddio n224__vddio 124.6e-3
ri963 n224__vddio n216__vddio 133e-3
ri964 n216__vddio n208__vddio 124.6e-3
ri965 n208__vddio n200__vddio 120e-3
ri966 n200__vddio n192__vddio 124.6e-3
ri967 n192__vddio n184__vddio 125.5e-3
ri968 n184__vddio n176__vddio 124.6e-3
ri969 n176__vddio n168__vddio 120e-3
ri970 n168__vddio n160__vddio 124.6e-3
ri971 n160__vddio n152__vddio 133e-3
ri972 n152__vddio n144__vddio 124.6e-3
ri973 n144__vddio n136__vddio 120e-3
ri974 n136__vddio n128__vddio 121.8e-3
ri975 n128__vddio n120__vddio 124.6e-3
ri976 n120__vddio n112__vddio 120e-3
ri977 n112__vddio n104__vddio 124.6e-3
ri978 n104__vddio n96__vddio 133e-3
ri979 n96__vddio n88__vddio 124.6e-3
ri980 n88__vddio n80__vddio 120e-3
ri981 n80__vddio n72__vddio 124.6e-3
ri982 n72__vddio n64__vddio 125.5e-3
ri983 n64__vddio n56__vddio 124.6e-3
ri984 n56__vddio n48__vddio 120e-3
ri985 n48__vddio n40__vddio 124.6e-3
ri986 n40__vddio n32__vddio 133e-3
ri987 n32__vddio n24__vddio 124.6e-3
ri988 n24__vddio n16__vddio 120e-3
ri989 n16__vddio n8__vddio 124.6e-3
ri990 n626__vddio n985__vddio 31.25e-3
ri991 n628__vddio n986__vddio 25e-3
ri992 n630__vddio n987__vddio 25e-3
ri993 n632__vddio n988__vddio 25e-3
rj1 n1__vss n2__vss 333.3e-3
rj2 n3__vss n4__vss 333.3e-3
rj3 n5__vss n6__vss 333.3e-3
rj4 n7__vss n8__vss 333.3e-3
rj5 n1__vddio n2__vddio 333.3e-3
rj6 n3__vddio n4__vddio 333.3e-3
rj7 n5__vddio n6__vddio 333.3e-3
rj8 n7__vddio n8__vddio 333.3e-3
rj9 n46__i18__net5 n47__i18__net5 1
rj10 n1__r_out n2__r_out 1
rj11 n3__r_out n4__r_out 1
rj12 n49__i18__net5 n48__i18__net5 500e-3
rj13 n9__vss n10__vss 333.3e-3
rj14 n11__vss n12__vss 333.3e-3
rj15 n13__vss n14__vss 333.3e-3
rj16 n15__vss n16__vss 333.3e-3
rj17 n9__vddio n10__vddio 333.3e-3
rj18 n11__vddio n12__vddio 333.3e-3
rj19 n13__vddio n14__vddio 333.3e-3
rj20 n15__vddio n16__vddio 333.3e-3
rj21 n56__i18__net5 n57__i18__net5 1
rj22 n17__r_out n23__r_out 1
rj23 n24__r_out n21__r_out 1
rj24 n59__i18__net5 n58__i18__net5 500e-3
rj25 n17__vss n18__vss 333.3e-3
rj26 n19__vss n20__vss 333.3e-3
rj27 n21__vss n22__vss 333.3e-3
rj28 n23__vss n24__vss 333.3e-3
rj29 n17__vddio n18__vddio 333.3e-3
rj30 n19__vddio n20__vddio 333.3e-3
rj31 n21__vddio n22__vddio 333.3e-3
rj32 n23__vddio n24__vddio 333.3e-3
rj33 n66__i18__net5 n67__i18__net5 1
rj34 n27__r_out n28__r_out 1
rj35 n29__r_out n30__r_out 1
rj36 n72__i18__net5 n71__i18__net5 500e-3
rj37 n25__vss n26__vss 333.3e-3
rj38 n27__vss n28__vss 333.3e-3
rj39 n29__vss n30__vss 333.3e-3
rj40 n31__vss n32__vss 333.3e-3
rj41 n25__vddio n26__vddio 333.3e-3
rj42 n27__vddio n28__vddio 333.3e-3
rj43 n29__vddio n30__vddio 333.3e-3
rj44 n31__vddio n32__vddio 333.3e-3
rj45 n76__i18__net5 n77__i18__net5 1
rj46 n40__r_out n41__r_out 1
rj47 n42__r_out n43__r_out 1
rj48 n82__i18__net5 n81__i18__net5 500e-3
rj49 n33__vss n34__vss 333.3e-3
rj50 n35__vss n36__vss 333.3e-3
rj51 n37__vss n38__vss 333.3e-3
rj52 n39__vss n40__vss 333.3e-3
rj53 n33__vddio n34__vddio 333.3e-3
rj54 n35__vddio n36__vddio 333.3e-3
rj55 n37__vddio n38__vddio 333.3e-3
rj56 n39__vddio n40__vddio 333.3e-3
rj57 n83__i18__net5 n84__i18__net5 500e-3
rj58 n53__r_out n54__r_out 1
rj59 n55__r_out n56__r_out 1
rj60 n89__i18__net5 n88__i18__net5 500e-3
rj61 n41__vss n42__vss 333.3e-3
rj62 n43__vss n44__vss 333.3e-3
rj63 n45__vss n46__vss 333.3e-3
rj64 n47__vss n48__vss 333.3e-3
rj65 n41__vddio n42__vddio 333.3e-3
rj66 n43__vddio n44__vddio 333.3e-3
rj67 n45__vddio n46__vddio 333.3e-3
rj68 n47__vddio n48__vddio 333.3e-3
rj69 n93__i18__net5 n94__i18__net5 1
rj70 n66__r_out n67__r_out 1
rj71 n68__r_out n69__r_out 1
rj72 n99__i18__net5 n98__i18__net5 500e-3
rj73 n49__vss n50__vss 333.3e-3
rj74 n51__vss n52__vss 333.3e-3
rj75 n53__vss n54__vss 333.3e-3
rj76 n55__vss n56__vss 333.3e-3
rj77 n49__vddio n50__vddio 333.3e-3
rj78 n51__vddio n52__vddio 333.3e-3
rj79 n53__vddio n54__vddio 333.3e-3
rj80 n55__vddio n56__vddio 333.3e-3
rj81 n106__i18__net5 n107__i18__net5 1
rj82 n82__r_out n88__r_out 1
rj83 n89__r_out n86__r_out 1
rj84 n108__i18__net5 n109__i18__net5 1
rj85 n57__vss n58__vss 333.3e-3
rj86 n59__vss n60__vss 333.3e-3
rj87 n61__vss n62__vss 333.3e-3
rj88 n63__vss n64__vss 333.3e-3
rj89 n57__vddio n58__vddio 333.3e-3
rj90 n59__vddio n60__vddio 333.3e-3
rj91 n61__vddio n62__vddio 333.3e-3
rj92 n63__vddio n64__vddio 333.3e-3
rj93 n113__i18__net5 n114__i18__net5 1
rj94 n92__r_out n93__r_out 1
rj95 n94__r_out n95__r_out 1
rj96 n118__i18__net5 n119__i18__net5 1
rj97 n65__vss n66__vss 333.3e-3
rj98 n67__vss n68__vss 333.3e-3
rj99 n69__vss n70__vss 333.3e-3
rj100 n71__vss n72__vss 333.3e-3
rj101 n65__vddio n66__vddio 333.3e-3
rj102 n67__vddio n68__vddio 333.3e-3
rj103 n69__vddio n70__vddio 333.3e-3
rj104 n71__vddio n72__vddio 333.3e-3
rj105 n126__i18__net5 n127__i18__net5 1
rj106 n105__r_out n106__r_out 1
rj107 n107__r_out n108__r_out 1
rj108 n132__i18__net5 n128__i18__net5 500e-3
rj109 n73__vss n74__vss 333.3e-3
rj110 n75__vss n76__vss 333.3e-3
rj111 n77__vss n78__vss 333.3e-3
rj112 n79__vss n80__vss 333.3e-3
rj113 n73__vddio n74__vddio 333.3e-3
rj114 n75__vddio n76__vddio 333.3e-3
rj115 n77__vddio n78__vddio 333.3e-3
rj116 n79__vddio n80__vddio 333.3e-3
rj117 n133__i18__net5 n134__i18__net5 1
rj118 n118__r_out n119__r_out 1
rj119 n120__r_out n121__r_out 1
rj120 n142__i18__net5 n141__i18__net5 500e-3
rj121 n81__vss n82__vss 333.3e-3
rj122 n83__vss n84__vss 333.3e-3
rj123 n85__vss n86__vss 333.3e-3
rj124 n87__vss n88__vss 333.3e-3
rj125 n81__vddio n82__vddio 333.3e-3
rj126 n83__vddio n84__vddio 333.3e-3
rj127 n85__vddio n86__vddio 333.3e-3
rj128 n87__vddio n88__vddio 333.3e-3
rj129 n146__i18__net5 n147__i18__net5 500e-3
rj130 n134__r_out n140__r_out 1
rj131 n141__r_out n138__r_out 1
rj132 n152__i18__net5 n151__i18__net5 500e-3
rj133 n89__vss n90__vss 333.3e-3
rj134 n91__vss n92__vss 333.3e-3
rj135 n93__vss n94__vss 333.3e-3
rj136 n95__vss n96__vss 333.3e-3
rj137 n89__vddio n90__vddio 333.3e-3
rj138 n91__vddio n92__vddio 333.3e-3
rj139 n93__vddio n94__vddio 333.3e-3
rj140 n95__vddio n96__vddio 333.3e-3
rj141 n156__i18__net5 n157__i18__net5 1
rj142 n147__r_out n153__r_out 1
rj143 n154__r_out n151__r_out 1
rj144 n159__i18__net5 n158__i18__net5 500e-3
rj145 n97__vss n98__vss 333.3e-3
rj146 n99__vss n100__vss 333.3e-3
rj147 n101__vss n102__vss 333.3e-3
rj148 n103__vss n104__vss 333.3e-3
rj149 n97__vddio n98__vddio 333.3e-3
rj150 n99__vddio n100__vddio 333.3e-3
rj151 n101__vddio n102__vddio 333.3e-3
rj152 n103__vddio n104__vddio 333.3e-3
rj153 n163__i18__net5 n167__i18__net5 500e-3
rj154 n157__r_out n158__r_out 1
rj155 n159__r_out n160__r_out 1
rj156 n169__i18__net5 n168__i18__net5 500e-3
rj157 n105__vss n106__vss 333.3e-3
rj158 n107__vss n108__vss 333.3e-3
rj159 n109__vss n110__vss 333.3e-3
rj160 n111__vss n112__vss 333.3e-3
rj161 n105__vddio n106__vddio 333.3e-3
rj162 n107__vddio n108__vddio 333.3e-3
rj163 n109__vddio n110__vddio 333.3e-3
rj164 n111__vddio n112__vddio 333.3e-3
rj165 n176__i18__net5 n177__i18__net5 1
rj166 n170__r_out n171__r_out 1
rj167 n172__r_out n173__r_out 1
rj168 n182__i18__net5 n178__i18__net5 500e-3
rj169 n113__vss n114__vss 333.3e-3
rj170 n115__vss n116__vss 333.3e-3
rj171 n117__vss n118__vss 333.3e-3
rj172 n119__vss n120__vss 333.3e-3
rj173 n113__vddio n114__vddio 333.3e-3
rj174 n115__vddio n116__vddio 333.3e-3
rj175 n117__vddio n118__vddio 333.3e-3
rj176 n119__vddio n120__vddio 333.3e-3
rj177 n183__i18__net5 n184__i18__net5 1
rj178 n183__r_out n184__r_out 1
rj179 n185__r_out n186__r_out 1
rj180 n192__i18__net5 n191__i18__net5 500e-3
rj181 n121__vss n122__vss 333.3e-3
rj182 n123__vss n124__vss 333.3e-3
rj183 n125__vss n126__vss 333.3e-3
rj184 n127__vss n128__vss 333.3e-3
rj185 n121__vddio n122__vddio 333.3e-3
rj186 n123__vddio n124__vddio 333.3e-3
rj187 n125__vddio n126__vddio 333.3e-3
rj188 n127__vddio n128__vddio 333.3e-3
rj189 n196__i18__net5 n197__i18__net5 1
rj190 n196__r_out n197__r_out 1
rj191 n198__r_out n199__r_out 1
rj192 n202__i18__net5 n198__i18__net5 500e-3
rj193 n129__vss n130__vss 333.3e-3
rj194 n131__vss n132__vss 333.3e-3
rj195 n133__vss n134__vss 333.3e-3
rj196 n135__vss n136__vss 333.3e-3
rj197 n129__vddio n130__vddio 333.3e-3
rj198 n131__vddio n132__vddio 333.3e-3
rj199 n133__vddio n134__vddio 333.3e-3
rj200 n135__vddio n136__vddio 333.3e-3
rj201 n206__i18__net5 n207__i18__net5 1
rj202 n212__r_out n218__r_out 1
rj203 n219__r_out n216__r_out 1
rj204 n212__i18__net5 n211__i18__net5 500e-3
rj205 n137__vss n138__vss 333.3e-3
rj206 n139__vss n140__vss 333.3e-3
rj207 n141__vss n142__vss 333.3e-3
rj208 n143__vss n144__vss 333.3e-3
rj209 n137__vddio n138__vddio 333.3e-3
rj210 n139__vddio n140__vddio 333.3e-3
rj211 n141__vddio n142__vddio 333.3e-3
rj212 n143__vddio n144__vddio 333.3e-3
rj213 n213__i18__net5 n217__i18__net5 500e-3
rj214 n222__r_out n223__r_out 1
rj215 n224__r_out n225__r_out 1
rj216 n222__i18__net5 n221__i18__net5 500e-3
rj217 n145__vss n146__vss 333.3e-3
rj218 n147__vss n148__vss 333.3e-3
rj219 n149__vss n150__vss 333.3e-3
rj220 n151__vss n152__vss 333.3e-3
rj221 n145__vddio n146__vddio 333.3e-3
rj222 n147__vddio n148__vddio 333.3e-3
rj223 n149__vddio n150__vddio 333.3e-3
rj224 n151__vddio n152__vddio 333.3e-3
rj225 n226__i18__net5 n227__i18__net5 1
rj226 n235__r_out n236__r_out 1
rj227 n237__r_out n238__r_out 1
rj228 n232__i18__net5 n231__i18__net5 500e-3
rj229 n153__vss n154__vss 333.3e-3
rj230 n155__vss n156__vss 333.3e-3
rj231 n157__vss n158__vss 333.3e-3
rj232 n159__vss n160__vss 333.3e-3
rj233 n153__vddio n154__vddio 333.3e-3
rj234 n155__vddio n156__vddio 333.3e-3
rj235 n157__vddio n158__vddio 333.3e-3
rj236 n159__vddio n160__vddio 333.3e-3
rj237 n233__i18__net5 n234__i18__net5 500e-3
rj238 n248__r_out n249__r_out 1
rj239 n250__r_out n251__r_out 1
rj240 n239__i18__net5 n238__i18__net5 500e-3
rj241 n161__vss n162__vss 333.3e-3
rj242 n163__vss n164__vss 333.3e-3
rj243 n165__vss n166__vss 333.3e-3
rj244 n167__vss n168__vss 333.3e-3
rj245 n161__vddio n162__vddio 333.3e-3
rj246 n163__vddio n164__vddio 333.3e-3
rj247 n165__vddio n166__vddio 333.3e-3
rj248 n167__vddio n168__vddio 333.3e-3
rj249 n243__i18__net5 n244__i18__net5 1
rj250 n261__r_out n262__r_out 1
rj251 n263__r_out n264__r_out 1
rj252 n249__i18__net5 n248__i18__net5 500e-3
rj253 n169__vss n170__vss 333.3e-3
rj254 n171__vss n172__vss 333.3e-3
rj255 n173__vss n174__vss 333.3e-3
rj256 n175__vss n176__vss 333.3e-3
rj257 n169__vddio n170__vddio 333.3e-3
rj258 n171__vddio n172__vddio 333.3e-3
rj259 n173__vddio n174__vddio 333.3e-3
rj260 n175__vddio n176__vddio 333.3e-3
rj261 n256__i18__net5 n257__i18__net5 1
rj262 n277__r_out n283__r_out 1
rj263 n284__r_out n281__r_out 1
rj264 n262__i18__net5 n261__i18__net5 500e-3
rj265 n177__vss n178__vss 333.3e-3
rj266 n179__vss n180__vss 333.3e-3
rj267 n181__vss n182__vss 333.3e-3
rj268 n183__vss n184__vss 333.3e-3
rj269 n177__vddio n178__vddio 333.3e-3
rj270 n179__vddio n180__vddio 333.3e-3
rj271 n181__vddio n182__vddio 333.3e-3
rj272 n183__vddio n184__vddio 333.3e-3
rj273 n263__i18__net5 n264__i18__net5 1
rj274 n287__r_out n288__r_out 1
rj275 n289__r_out n290__r_out 1
rj276 n272__i18__net5 n271__i18__net5 500e-3
rj277 n185__vss n186__vss 333.3e-3
rj278 n187__vss n188__vss 333.3e-3
rj279 n189__vss n190__vss 333.3e-3
rj280 n191__vss n192__vss 333.3e-3
rj281 n185__vddio n186__vddio 333.3e-3
rj282 n187__vddio n188__vddio 333.3e-3
rj283 n189__vddio n190__vddio 333.3e-3
rj284 n191__vddio n192__vddio 333.3e-3
rj285 n273__i18__net5 n274__i18__net5 1
rj286 n300__r_out n301__r_out 1
rj287 n302__r_out n303__r_out 1
rj288 n282__i18__net5 n281__i18__net5 500e-3
rj289 n193__vss n194__vss 333.3e-3
rj290 n195__vss n196__vss 333.3e-3
rj291 n197__vss n198__vss 333.3e-3
rj292 n199__vss n200__vss 333.3e-3
rj293 n193__vddio n194__vddio 333.3e-3
rj294 n195__vddio n196__vddio 333.3e-3
rj295 n197__vddio n198__vddio 333.3e-3
rj296 n199__vddio n200__vddio 333.3e-3
rj297 n286__i18__net5 n287__i18__net5 1
rj298 n313__r_out n314__r_out 1
rj299 n315__r_out n316__r_out 1
rj300 n292__i18__net5 n291__i18__net5 500e-3
rj301 n201__vss n202__vss 333.3e-3
rj302 n203__vss n204__vss 333.3e-3
rj303 n205__vss n206__vss 333.3e-3
rj304 n207__vss n208__vss 333.3e-3
rj305 n201__vddio n202__vddio 333.3e-3
rj306 n203__vddio n204__vddio 333.3e-3
rj307 n205__vddio n206__vddio 333.3e-3
rj308 n207__vddio n208__vddio 333.3e-3
rj309 n296__i18__net5 n297__i18__net5 1
rj310 n326__r_out n327__r_out 1
rj311 n328__r_out n329__r_out 1
rj312 n302__i18__net5 n301__i18__net5 500e-3
rj313 n209__vss n210__vss 333.3e-3
rj314 n211__vss n212__vss 333.3e-3
rj315 n213__vss n214__vss 333.3e-3
rj316 n215__vss n216__vss 333.3e-3
rj317 n209__vddio n210__vddio 333.3e-3
rj318 n211__vddio n212__vddio 333.3e-3
rj319 n213__vddio n214__vddio 333.3e-3
rj320 n215__vddio n216__vddio 333.3e-3
rj321 n306__i18__net5 n307__i18__net5 1
rj322 n342__r_out n348__r_out 1
rj323 n349__r_out n346__r_out 1
rj324 n309__i18__net5 n308__i18__net5 500e-3
rj325 n217__vss n218__vss 333.3e-3
rj326 n219__vss n220__vss 333.3e-3
rj327 n221__vss n222__vss 333.3e-3
rj328 n223__vss n224__vss 333.3e-3
rj329 n217__vddio n218__vddio 333.3e-3
rj330 n219__vddio n220__vddio 333.3e-3
rj331 n221__vddio n222__vddio 333.3e-3
rj332 n223__vddio n224__vddio 333.3e-3
rj333 n316__i18__net5 n317__i18__net5 1
rj334 n352__r_out n353__r_out 1
rj335 n354__r_out n355__r_out 1
rj336 n319__i18__net5 n318__i18__net5 500e-3
rj337 n225__vss n226__vss 333.3e-3
rj338 n227__vss n228__vss 333.3e-3
rj339 n229__vss n230__vss 333.3e-3
rj340 n231__vss n232__vss 333.3e-3
rj341 n225__vddio n226__vddio 333.3e-3
rj342 n227__vddio n228__vddio 333.3e-3
rj343 n229__vddio n230__vddio 333.3e-3
rj344 n231__vddio n232__vddio 333.3e-3
rj345 n323__i18__net5 n324__i18__net5 1
rj346 n365__r_out n366__r_out 1
rj347 n367__r_out n368__r_out 1
rj348 n332__i18__net5 n331__i18__net5 500e-3
rj349 n233__vss n234__vss 333.3e-3
rj350 n235__vss n236__vss 333.3e-3
rj351 n237__vss n238__vss 333.3e-3
rj352 n239__vss n240__vss 333.3e-3
rj353 n233__vddio n234__vddio 333.3e-3
rj354 n235__vddio n236__vddio 333.3e-3
rj355 n237__vddio n238__vddio 333.3e-3
rj356 n239__vddio n240__vddio 333.3e-3
rj357 n333__i18__net5 n334__i18__net5 1
rj358 n378__r_out n379__r_out 1
rj359 n380__r_out n381__r_out 1
rj360 n342__i18__net5 n341__i18__net5 500e-3
rj361 n241__vss n242__vss 333.3e-3
rj362 n243__vss n244__vss 333.3e-3
rj363 n245__vss n246__vss 333.3e-3
rj364 n247__vss n248__vss 333.3e-3
rj365 n241__vddio n242__vddio 333.3e-3
rj366 n243__vddio n244__vddio 333.3e-3
rj367 n245__vddio n246__vddio 333.3e-3
rj368 n247__vddio n248__vddio 333.3e-3
rj369 n343__i18__net5 n344__i18__net5 1
rj370 n391__r_out n392__r_out 1
rj371 n393__r_out n394__r_out 1
rj372 n352__i18__net5 n351__i18__net5 500e-3
rj373 n249__vss n250__vss 333.3e-3
rj374 n251__vss n252__vss 333.3e-3
rj375 n253__vss n254__vss 333.3e-3
rj376 n255__vss n256__vss 333.3e-3
rj377 n249__vddio n250__vddio 333.3e-3
rj378 n251__vddio n252__vddio 333.3e-3
rj379 n253__vddio n254__vddio 333.3e-3
rj380 n255__vddio n256__vddio 333.3e-3
rj381 n353__i18__net5 n354__i18__net5 1
rj382 n407__r_out n413__r_out 1
rj383 n414__r_out n411__r_out 1
rj384 n359__i18__net5 n358__i18__net5 500e-3
rj385 n257__vss n258__vss 333.3e-3
rj386 n259__vss n260__vss 333.3e-3
rj387 n261__vss n262__vss 333.3e-3
rj388 n263__vss n264__vss 333.3e-3
rj389 n257__vddio n258__vddio 333.3e-3
rj390 n259__vddio n260__vddio 333.3e-3
rj391 n261__vddio n262__vddio 333.3e-3
rj392 n263__vddio n264__vddio 333.3e-3
rj393 n363__i18__net5 n364__i18__net5 1
rj394 n420__r_out n426__r_out 1
rj395 n427__r_out n424__r_out 1
rj396 n372__i18__net5 n371__i18__net5 500e-3
rj397 n265__vss n266__vss 333.3e-3
rj398 n267__vss n268__vss 333.3e-3
rj399 n269__vss n270__vss 333.3e-3
rj400 n271__vss n272__vss 333.3e-3
rj401 n265__vddio n266__vddio 333.3e-3
rj402 n267__vddio n268__vddio 333.3e-3
rj403 n269__vddio n270__vddio 333.3e-3
rj404 n271__vddio n272__vddio 333.3e-3
rj405 n373__i18__net5 n374__i18__net5 500e-3
rj406 n432__r_out n433__r_out 1
rj407 n434__r_out n435__r_out 1
rj408 n382__i18__net5 n381__i18__net5 500e-3
rj409 n273__vss n274__vss 333.3e-3
rj410 n275__vss n276__vss 333.3e-3
rj411 n277__vss n278__vss 333.3e-3
rj412 n279__vss n280__vss 333.3e-3
rj413 n273__vddio n274__vddio 333.3e-3
rj414 n275__vddio n276__vddio 333.3e-3
rj415 n277__vddio n278__vddio 333.3e-3
rj416 n279__vddio n280__vddio 333.3e-3
rj417 n383__i18__net5 n384__i18__net5 500e-3
rj418 n448__r_out n454__r_out 1
rj419 n455__r_out n452__r_out 1
rj420 n389__i18__net5 n388__i18__net5 500e-3
rj421 n281__vss n282__vss 333.3e-3
rj422 n283__vss n284__vss 333.3e-3
rj423 n285__vss n286__vss 333.3e-3
rj424 n287__vss n288__vss 333.3e-3
rj425 n281__vddio n282__vddio 333.3e-3
rj426 n283__vddio n284__vddio 333.3e-3
rj427 n285__vddio n286__vddio 333.3e-3
rj428 n287__vddio n288__vddio 333.3e-3
rj429 n393__i18__net5 n394__i18__net5 500e-3
rj430 n464__r_out n470__r_out 1
rj431 n471__r_out n468__r_out 1
rj432 n401__i18__net5 n402__i18__net5 1
rj433 n289__vss n290__vss 333.3e-3
rj434 n291__vss n292__vss 333.3e-3
rj435 n293__vss n294__vss 333.3e-3
rj436 n295__vss n296__vss 333.3e-3
rj437 n289__vddio n290__vddio 333.3e-3
rj438 n291__vddio n292__vddio 333.3e-3
rj439 n293__vddio n294__vddio 333.3e-3
rj440 n295__vddio n296__vddio 333.3e-3
rj441 n403__i18__net5 n404__i18__net5 1
rj442 n474__r_out n475__r_out 1
rj443 n476__r_out n477__r_out 1
rj444 n412__i18__net5 n411__i18__net5 500e-3
rj445 n297__vss n298__vss 333.3e-3
rj446 n299__vss n300__vss 333.3e-3
rj447 n301__vss n302__vss 333.3e-3
rj448 n303__vss n304__vss 333.3e-3
rj449 n297__vddio n298__vddio 333.3e-3
rj450 n299__vddio n300__vddio 333.3e-3
rj451 n301__vddio n302__vddio 333.3e-3
rj452 n303__vddio n304__vddio 333.3e-3
rj453 n416__i18__net5 n417__i18__net5 1
rj454 n487__r_out n488__r_out 1
rj455 n489__r_out n490__r_out 1
rj456 n422__i18__net5 n418__i18__net5 500e-3
rj457 n305__vss n306__vss 333.3e-3
rj458 n307__vss n308__vss 333.3e-3
rj459 n309__vss n310__vss 333.3e-3
rj460 n311__vss n312__vss 333.3e-3
rj461 n305__vddio n306__vddio 333.3e-3
rj462 n307__vddio n308__vddio 333.3e-3
rj463 n309__vddio n310__vddio 333.3e-3
rj464 n311__vddio n312__vddio 333.3e-3
rj465 n2__x3 n4__x3 1
rj466 n4__x2 n2__x2 1
rj467 n2__x1 n4__x1 1
rj468 n4__x0 n2__x0 1
rj469 n426__i18__net5 n427__i18__net5 500e-3
rj470 n500__r_out n501__r_out 1
rj471 n502__r_out n503__r_out 1
rj472 n9__i14__i17__net1 n6__i14__i17__net1 560.4e-3
rj473 n5__i14__i17__net8 n2__i14__i17__net8 560.4e-3
rj474 n431__i18__net5 n432__i18__net5 500e-3
rj475 n313__vss n314__vss 333.3e-3
rj476 n315__vss n316__vss 333.3e-3
rj477 n317__vss n318__vss 333.3e-3
rj478 n319__vss n320__vss 333.3e-3
rj479 n313__vddio n314__vddio 333.3e-3
rj480 n315__vddio n316__vddio 333.3e-3
rj481 n317__vddio n318__vddio 333.3e-3
rj482 n319__vddio n320__vddio 333.3e-3
rj484 n21__i14__net9 n17__i14__net9 479.5e-3
rj486 n23__i14__net9 n18__i14__net9 479.5e-3
rj488 n25__i14__net9 n19__i14__net9 479.5e-3
rj490 n27__i14__net9 n20__i14__net9 479.5e-3
rj491 n433__i18__net5 n434__i18__net5 1
rj493 n37__i14__net10 n18__i14__net10 1.0681
rj495 n39__i14__net10 n22__i14__net10 1.0681
rj497 n41__i14__net10 n24__i14__net10 1.0681
rj499 n43__i14__net10 n28__i14__net10 1.0681
rj500 n513__r_out n514__r_out 1
rj501 n515__r_out n516__r_out 1
rj502 n438__i18__net5 n439__i18__net5 500e-3
rj503 n18__i14__i17__net1 n13__i14__i17__net1 932.5e-3
rj504 n13__i14__i17__net1 n10__i14__i17__net1 46.98e-3
rj505 n9__i14__i17__net3 n8__i14__i17__net3 979.5e-3
rj506 n8__i14__i17__net3 n6__i14__i17__net3 719.8e-3
rj507 n321__vss n322__vss 333.3e-3
rj508 n323__vss n324__vss 333.3e-3
rj509 n325__vss n326__vss 333.3e-3
rj510 n327__vss n328__vss 333.3e-3
rj511 n321__vddio n322__vddio 333.3e-3
rj512 n323__vddio n324__vddio 333.3e-3
rj513 n325__vddio n326__vddio 333.3e-3
rj514 n327__vddio n328__vddio 333.3e-3
rj515 n9__i14__net3 n10__i14__net3 1
rj516 n11__i14__net3 n12__i14__net3 1
rj517 n13__i14__net3 n14__i14__net3 1
rj518 n15__i14__net3 n16__i14__net3 1
rj519 n10__i14__i17__net7 n8__i14__i17__net7 374.8e-3
rj520 n8__i14__i17__net7 n7__i14__i17__net7 693.3e-3
rj522 n16__ck n18__ck 568.1e-3
rj523 n18__ck n8__ck 826.1e-3
rj524 n13__ck n18__ck 500e-3
rj525 n446__i18__net5 n447__i18__net5 1
rj526 n16__i14__i13__net1 n14__i14__i13__net1 669.1e-3
rj527 n14__i14__i13__net1 n11__i14__i13__net1 1.1446
rj528 n16__i14__i16__net1 n14__i14__i16__net1 669.1e-3
rj529 n14__i14__i16__net1 n11__i14__i16__net1 1.1446
rj530 n16__i14__i10__net1 n14__i14__i10__net1 669.1e-3
rj531 n14__i14__i10__net1 n11__i14__i10__net1 1.1446
rj532 n16__i14__i9__net1 n14__i14__i9__net1 669.1e-3
rj533 n14__i14__i9__net1 n11__i14__i9__net1 1.1446
rj534 n535__r_out n529__r_out 1
rj535 n533__r_out n536__r_out 1
rj537 n22__reset n14__reset 1.1072
rj538 n17__reset n22__reset 500e-3
rj539 n19__reset n15__reset 1.6025
rj540 n15__reset n24__reset 75.39e-3
rj541 n24__reset n12__reset 4.832e-3
rj542 n8__reset n24__reset 500e-3
rj543 n448__i18__net5 n449__i18__net5 1
rj544 n5__i14__i13__net2 n4__i14__i13__net2 1.2876
rj545 n5__i14__i16__net2 n4__i14__i16__net2 1.2876
rj546 n5__i14__i10__net2 n4__i14__i10__net2 1.2876
rj547 n5__i14__i9__net2 n4__i14__i9__net2 1.2876
rj548 n329__vss n330__vss 333.3e-3
rj549 n331__vss n332__vss 333.3e-3
rj550 n333__vss n334__vss 333.3e-3
rj551 n335__vss n336__vss 333.3e-3
rj552 n329__vddio n330__vddio 333.3e-3
rj553 n331__vddio n332__vddio 333.3e-3
rj554 n333__vddio n334__vddio 333.3e-3
rj555 n335__vddio n336__vddio 333.3e-3
rj556 n16__i14__i17__i2__net1 n14__i14__i17__i2__net1 669.1e-3
rj557 n14__i14__i17__i2__net1 n11__i14__i17__i2__net1 1.1446
rj558 n16__i14__i17__i3__net1 n14__i14__i17__i3__net1 669.1e-3
rj559 n14__i14__i17__i3__net1 n11__i14__i17__i3__net1 1.1446
rj560 n456__i18__net5 n457__i18__net5 1
rj561 n5__i14__i17__i2__net2 n4__i14__i17__i2__net2 1.2876
rj562 n5__i14__i17__i3__net2 n4__i14__i17__i3__net2 1.2876
rj563 n548__r_out n542__r_out 1
rj564 n546__r_out n549__r_out 1
rj565 n45__i14__net9 n41__i14__net9 731.9e-3
rj566 n46__i14__net9 n42__i14__net9 731.9e-3
rj567 n47__i14__net9 n43__i14__net9 731.9e-3
rj568 n48__i14__net9 n44__i14__net9 731.9e-3
rj569 n53__i14__net10 n49__i14__net10 829e-3
rj570 n54__i14__net10 n50__i14__net10 829e-3
rj571 n55__i14__net10 n51__i14__net10 829e-3
rj572 n56__i14__net10 n52__i14__net10 829e-3
rj573 n461__i18__net5 n462__i18__net5 500e-3
rj574 n337__vss n338__vss 333.3e-3
rj575 n339__vss n340__vss 333.3e-3
rj576 n341__vss n342__vss 333.3e-3
rj577 n343__vss n344__vss 333.3e-3
rj578 n337__vddio n338__vddio 333.3e-3
rj579 n339__vddio n340__vddio 333.3e-3
rj580 n341__vddio n342__vddio 333.3e-3
rj581 n343__vddio n344__vddio 333.3e-3
rj582 n466__i18__net5 n467__i18__net5 1
rj583 n11__i14__i17__net3 n10__i14__i17__net3 731.9e-3
rj584 n20__i14__i17__net1 n19__i14__i17__net1 731.9e-3
rj585 n21__ck n15__ck 829e-3
rj586 n12__i14__i17__net7 n11__i14__i17__net7 829e-3
rj587 n561__r_out n555__r_out 1
rj588 n559__r_out n562__r_out 1
rj589 n1__vdd n2__vdd 166.7e-3
rj590 n3__vdd n4__vdd 166.7e-3
rj591 n5__vdd n6__vdd 166.7e-3
rj592 n468__i18__net5 n469__i18__net5 500e-3
rj593 n345__vss n346__vss 333.3e-3
rj594 n347__vss n348__vss 333.3e-3
rj595 n349__vss n350__vss 333.3e-3
rj596 n351__vss n352__vss 333.3e-3
rj597 n345__vddio n346__vddio 333.3e-3
rj598 n347__vddio n348__vddio 333.3e-3
rj599 n349__vddio n350__vddio 333.3e-3
rj600 n351__vddio n352__vddio 333.3e-3
rj601 n17__i14__net4 n10__i14__net4 631.1e-3
rj602 n18__i14__net4 n11__i14__net4 631.1e-3
rj603 n19__i14__net4 n14__i14__net4 631.1e-3
rj604 n20__i14__net4 n15__i14__net4 631.1e-3
rj605 n473__i18__net5 n474__i18__net5 500e-3
rj606 n14__i14__i13__net5 n11__i14__i13__net5 1.447
rj607 n14__i14__i16__net5 n11__i14__i16__net5 1.447
rj608 n14__i14__i10__net5 n11__i14__i10__net5 1.447
rj609 n14__i14__i9__net5 n11__i14__i9__net5 1.447
rj610 n574__r_out n568__r_out 1
rj611 n572__r_out n575__r_out 1
rj612 n475__i18__net5 n476__i18__net5 500e-3
rj613 n10__i14__i17__net6 n8__i14__i17__net6 2.7224
rj614 n11__i14__i17__net6 n9__i14__i17__net6 2.723
rj615 n9__i14__i17__net6 n6__i14__i17__net6 555.3e-3
rj616 n12__i14__i13__net4 n7__i14__i13__net4 524.3e-3
rj617 n12__i14__i16__net4 n7__i14__i16__net4 524.3e-3
rj618 n12__i14__i10__net4 n7__i14__i10__net4 524.3e-3
rj619 n12__i14__i9__net4 n7__i14__i9__net4 524.3e-3
rj620 n353__vss n354__vss 333.3e-3
rj621 n355__vss n356__vss 333.3e-3
rj622 n357__vss n358__vss 333.3e-3
rj623 n359__vss n360__vss 333.3e-3
rj624 n353__vddio n354__vddio 333.3e-3
rj625 n355__vddio n356__vddio 333.3e-3
rj626 n357__vddio n358__vddio 333.3e-3
rj627 n359__vddio n360__vddio 333.3e-3
rj628 n14__i14__i17__i2__net5 n11__i14__i17__i2__net5 1.447
rj629 n14__i14__i17__i3__net5 n11__i14__i17__i3__net5 1.447
rj630 n477__i18__net5 n478__i18__net5 500e-3
rj631 n581__r_out n588__r_out 500e-3
rj632 n589__r_out n585__r_out 500e-3
rj633 n13__i14__i13__net4 n9__i14__i13__net4 712.6e-3
rj634 n13__i14__i16__net4 n9__i14__i16__net4 712.6e-3
rj635 n13__i14__i10__net4 n9__i14__i10__net4 712.6e-3
rj636 n13__i14__i9__net4 n9__i14__i9__net4 712.6e-3
rj637 n12__i14__i17__i2__net4 n7__i14__i17__i2__net4 524.3e-3
rj638 n12__i14__i17__i3__net4 n7__i14__i17__i3__net4 524.3e-3
rj639 n479__i18__net5 n480__i18__net5 500e-3
rj640 n361__vss n362__vss 333.3e-3
rj641 n363__vss n364__vss 333.3e-3
rj642 n365__vss n366__vss 333.3e-3
rj643 n367__vss n368__vss 333.3e-3
rj644 n361__vddio n362__vddio 333.3e-3
rj645 n363__vddio n364__vddio 333.3e-3
rj646 n365__vddio n366__vddio 333.3e-3
rj647 n367__vddio n368__vddio 333.3e-3
rj648 n481__i18__net5 n482__i18__net5 1
rj649 n13__i14__i17__i2__net4 n9__i14__i17__i2__net4 1.2126
rj650 n13__i14__i17__i3__net4 n9__i14__i17__i3__net4 1.2126
rj651 n600__r_out n594__r_out 1
rj652 n598__r_out n601__r_out 1
rj653 n17__i14__i17__net8 n4__i14__i17__net8 3.0703
rj654 n4__x_out_3 n2__x_out_3 1
rj655 n2__x_out_2 n4__x_out_2 1
rj656 n4__x_out_1 n2__x_out_1 1
rj657 n2__x_out_0 n4__x_out_0 1
rj662 n23__i14__i17__net1 n8__i14__i17__net1 3.077
rj663 n484__i18__net5 n483__i18__net5 500e-3
rj664 n369__vss n370__vss 333.3e-3
rj665 n371__vss n372__vss 333.3e-3
rj666 n373__vss n374__vss 333.3e-3
rj667 n375__vss n376__vss 333.3e-3
rj668 n369__vddio n370__vddio 333.3e-3
rj669 n371__vddio n372__vddio 333.3e-3
rj670 n373__vddio n374__vddio 333.3e-3
rj671 n375__vddio n376__vddio 333.3e-3
rj672 n5__y3 n2__y3 500e-3
rj673 n2__y2 n4__y2 500e-3
rj674 n5__y1 n2__y1 500e-3
rj675 n2__y0 n4__y0 500e-3
rj676 n485__i18__net5 n486__i18__net5 500e-3
rj677 n15__i14__i17__net7 n18__i14__i17__net7 500e-3
rj678 n11__i14__i17__net11 n9__i14__i17__net11 500e-3
rj680 n31__i14__i17__net1 n24__i14__i17__net1 500e-3
rj681 n27__i14__i17__net1 n31__i14__i17__net1 500e-3
rj682 n607__r_out n613__r_out 1
rj683 n614__r_out n611__r_out 1
rj684 n487__i18__net5 n488__i18__net5 1
rj685 n8__i14__i17__net10 n9__i14__i17__net10 1
rj686 n377__vss n378__vss 333.3e-3
rj687 n379__vss n380__vss 333.3e-3
rj688 n381__vss n382__vss 333.3e-3
rj689 n383__vss n384__vss 333.3e-3
rj690 n377__vddio n378__vddio 333.3e-3
rj691 n379__vddio n380__vddio 333.3e-3
rj692 n381__vddio n382__vddio 333.3e-3
rj693 n383__vddio n384__vddio 333.3e-3
rj694 n489__i18__net5 n490__i18__net5 500e-3
rj696 n61__i14__net9 n57__i14__net9 479.5e-3
rj698 n63__i14__net9 n58__i14__net9 479.5e-3
rj700 n65__i14__net9 n59__i14__net9 479.5e-3
rj702 n67__i14__net9 n60__i14__net9 479.5e-3
rj703 n12__i14__i17__net9 n11__i14__i17__net9 1
rj704 n626__r_out n620__r_out 1
rj705 n624__r_out n627__r_out 1
rj707 n78__i14__net10 n66__i14__net10 1.0681
rj709 n79__i14__net10 n70__i14__net10 1.0681
rj711 n82__i14__net10 n72__i14__net10 1.0681
rj713 n83__i14__net10 n76__i14__net10 1.0681
rj714 n491__i18__net5 n492__i18__net5 500e-3
rj715 n385__vss n386__vss 333.3e-3
rj716 n387__vss n388__vss 333.3e-3
rj717 n389__vss n390__vss 333.3e-3
rj718 n391__vss n392__vss 333.3e-3
rj719 n385__vddio n386__vddio 333.3e-3
rj720 n387__vddio n388__vddio 333.3e-3
rj721 n389__vddio n390__vddio 333.3e-3
rj722 n391__vddio n392__vddio 333.3e-3
rj723 n493__i18__net5 n494__i18__net5 500e-3
rj724 n38__i14__net3 n49__i14__net3 1
rj725 n50__i14__net3 n40__i14__net3 1
rj726 n44__i14__net3 n51__i14__net3 1
rj727 n52__i14__net3 n46__i14__net3 1
rj728 n16__i14__i11__net1 n14__i14__i11__net1 669.1e-3
rj729 n14__i14__i11__net1 n11__i14__i11__net1 1.1446
rj730 n16__i14__i14__net1 n14__i14__i14__net1 669.1e-3
rj731 n14__i14__i14__net1 n11__i14__i14__net1 1.1446
rj732 n16__i14__i15__net1 n14__i14__i15__net1 669.1e-3
rj733 n14__i14__i15__net1 n11__i14__i15__net1 1.1446
rj734 n16__i14__i12__net1 n14__i14__i12__net1 669.1e-3
rj735 n14__i14__i12__net1 n11__i14__i12__net1 1.1446
rj736 n639__r_out n633__r_out 1
rj737 n637__r_out n640__r_out 1
rj738 n495__i18__net5 n496__i18__net5 1
rj739 n5__i14__i11__net2 n4__i14__i11__net2 1.2876
rj740 n5__i14__i14__net2 n4__i14__i14__net2 1.2876
rj741 n5__i14__i15__net2 n4__i14__i15__net2 1.2876
rj742 n5__i14__i12__net2 n4__i14__i12__net2 1.2876
rj743 n393__vss n394__vss 333.3e-3
rj744 n395__vss n396__vss 333.3e-3
rj745 n397__vss n398__vss 333.3e-3
rj746 n399__vss n400__vss 333.3e-3
rj747 n393__vddio n394__vddio 333.3e-3
rj748 n395__vddio n396__vddio 333.3e-3
rj749 n397__vddio n398__vddio 333.3e-3
rj750 n399__vddio n400__vddio 333.3e-3
rj751 n401__vss n402__vss 166.7e-3
rj752 n403__vss n404__vss 166.7e-3
rj753 n405__vss n406__vss 166.7e-3
rj754 n407__vss n408__vss 166.7e-3
rj755 n49__reset n48__reset 201.9e-3
rj756 n48__reset n46__reset 196.4e-3
rj757 n25__i14__i17__net8 n24__i14__i17__net8 1.1242
rj758 n24__i14__i17__net8 n26__i14__i17__net8 234.3e-3
rj759 n26__i14__i17__net8 n27__i14__i17__net8 433.7e-3
rj760 n26__i14__i17__net8 n23__i14__i17__net8 39.53e-3
rj761 n27__i14__i17__net8 n18__i14__i17__net8 9.367e-3
rj762 n21__i14__i17__net8 n27__i14__i17__net8 500e-3
rj763 n497__i18__net5 n498__i18__net5 1
rj764 n15__i14__i17__net11 n16__i14__i17__net11 755.3e-3
rj765 n16__i14__i17__net11 n17__i14__i17__net11 594.4e-3
rj766 n17__i14__i17__net11 n8__i14__i17__net11 282.4e-3
rj767 n16__i14__i17__net11 n14__i14__i17__net11 40.26e-3
rj768 n17__i14__i17__net11 n13__i14__i17__net11 513.3e-3
rj769 n652__r_out n646__r_out 1
rj770 n650__r_out n653__r_out 1
rj771 n19__i14__i17__net10 n21__i14__i17__net10 760.8e-3
rj772 n21__i14__i17__net10 n22__i14__i17__net10 206e-3
rj773 n22__i14__i17__net10 n10__i14__i17__net10 449.9e-3
rj774 n17__i14__i17__net10 n21__i14__i17__net10 500e-3
rj775 n12__i14__i17__net10 n22__i14__i17__net10 500e-3
rj776 n19__i14__i17__net9 n21__i14__i17__net9 700.8e-3
rj777 n21__i14__i17__net9 n13__i14__i17__net9 100.8e-3
rj778 n13__i14__i17__net9 n9__i14__i17__net9 648.2e-3
rj779 n14__i14__i17__net9 n21__i14__i17__net9 500e-3
rj780 n499__i18__net5 n500__i18__net5 125e-3
rj781 n77__i14__net9 n73__i14__net9 731.9e-3
rj782 n78__i14__net9 n74__i14__net9 731.9e-3
rj783 n79__i14__net9 n75__i14__net9 731.9e-3
rj784 n80__i14__net9 n76__i14__net9 731.9e-3
rj785 n93__i14__net10 n77__i14__net10 829e-3
rj786 n94__i14__net10 n80__i14__net10 829e-3
rj787 n95__i14__net10 n81__i14__net10 829e-3
rj788 n96__i14__net10 n84__i14__net10 829e-3
rj789 n417__vss n418__vss 333.3e-3
rj790 n419__vss n420__vss 333.3e-3
rj791 n421__vss n422__vss 333.3e-3
rj792 n423__vss n424__vss 333.3e-3
rj793 n401__vddio n402__vddio 333.3e-3
rj794 n403__vddio n404__vddio 333.3e-3
rj795 n405__vddio n406__vddio 333.3e-3
rj796 n407__vddio n408__vddio 333.3e-3
rj797 n58__i14__net4 n59__i14__net4 761.7e-3
rj798 n59__i14__net4 n60__i14__net4 195.5e-3
rj799 n60__i14__net4 n50__i14__net4 694.1e-3
rj800 n56__i14__net4 n59__i14__net4 500e-3
rj801 n53__i14__net4 n60__i14__net4 500e-3
rj802 n29__i14__net7 n28__i14__net7 1.4113
rj804 n33__i14__net7 n32__i14__net7 500e-3
rj805 n31__i14__net11 n30__i14__net11 703.9e-3
rj806 n30__i14__net11 n28__i14__net11 1.1776
rj808 n71__i14__net4 n70__i14__net4 201.8e-3
rj809 n70__i14__net4 n61__i14__net4 586.8e-3
rj814 n417__vddio n418__vddio 166.7e-3
rj815 n433__vss n434__vss 166.7e-3
rj820 n68__i14__net3 n63__i14__net3 652.6e-3
rj821 n63__i14__net3 n69__i14__net3 30.34e-3
rj822 n69__i14__net3 n58__i14__net3 696.5e-3
rj823 n61__i14__net3 n69__i14__net3 500e-3
rj824 n72__i14__net4 n62__i14__net4 1.4221
rj825 n73__i14__net4 n64__i14__net4 1.4221
rj826 n74__i14__net4 n66__i14__net4 1.4221
rj827 n75__i14__net4 n69__i14__net4 922.1e-3
rj828 n14__i14__i11__net5 n11__i14__i11__net5 1.447
rj829 n14__i14__i14__net5 n11__i14__i14__net5 1.447
rj830 n14__i14__i15__net5 n11__i14__i15__net5 1.447
rj831 n14__i14__i12__net5 n11__i14__i12__net5 1.447
rj832 n8__i14__i11__net4 n7__i14__i11__net4 1.0243
rj833 n8__i14__i14__net4 n7__i14__i14__net4 1.0243
rj834 n8__i14__i15__net4 n7__i14__i15__net4 1.0243
rj835 n8__i14__i12__net4 n7__i14__i12__net4 1.0243
rj836 n429__vddio n430__vddio 333.3e-3
rj837 n431__vddio n432__vddio 333.3e-3
rj838 n433__vddio n434__vddio 333.3e-3
rj839 n43__i18__net4 n44__i18__net4 1
rj840 n34__i14__net7 n35__i14__net7 1
rj841 n33__i14__net11 n34__i14__net11 1
rj842 n502__i18__net5 n503__i18__net5 1
rj843 n504__i18__net5 n505__i18__net5 1
rj844 n13__i14__i11__net4 n10__i14__i11__net4 1.2126
rj845 n13__i14__i14__net4 n10__i14__i14__net4 1.2126
rj846 n13__i14__i15__net4 n10__i14__i15__net4 1.2126
rj847 n13__i14__i12__net4 n10__i14__i12__net4 1.2126
rj848 n51__i18__net4 n52__i18__net4 500e-3
rj849 n451__vddio n452__vddio 333.3e-3
rj850 n453__vddio n454__vddio 333.3e-3
rj851 n455__vddio n456__vddio 333.3e-3
rj852 n38__i14__net7 n37__i14__net7 500e-3
rj853 n36__i14__net11 n37__i14__net11 500e-3
rj854 n56__i18__net4 n57__i18__net4 500e-3
rj855 n81__i14__net9 n95__i14__net9 239.6e-3
rj856 n95__i14__net9 n96__i14__net9 200.8e-3
rj857 n96__i14__net9 n93__i14__net9 698.6e-3
rj858 n87__i14__net9 n95__i14__net9 500e-3
rj859 n90__i14__net9 n96__i14__net9 500e-3
rj860 n524__i18__net5 n518__i18__net5 1
rj861 n522__i18__net5 n525__i18__net5 1
rj862 n106__i14__net10 n107__i14__net10 575.7e-3
rj863 n107__i14__net10 n108__i14__net10 200.8e-3
rj864 n108__i14__net10 n98__i14__net10 698.6e-3
rj865 n104__i14__net10 n107__i14__net10 500e-3
rj866 n101__i14__net10 n108__i14__net10 500e-3
rj867 n8__y_out_3 n6__y_out_3 594.2e-3
rj868 n8__y_out_2 n5__y_out_2 594.2e-3
rj869 n8__y_out_1 n6__y_out_1 594.2e-3
rj870 n10__y_out_0 n7__y_out_0 594.2e-3
rj875 n58__i18__net4 n62__i18__net4 500e-3
rj876 n5__ck4 n4__ck4 1.2707
rj877 n457__vddio n458__vddio 333.3e-3
rj878 n459__vddio n460__vddio 333.3e-3
rj879 n461__vddio n462__vddio 333.3e-3
rj880 n66__i18__net4 n67__i18__net4 1
rj881 n537__i18__net5 n531__i18__net5 1
rj882 n535__i18__net5 n538__i18__net5 1
rj883 n17__x_out_2 n18__x_out_2 646.3e-3
rj884 n18__x_out_2 n14__x_out_2 24.35e-3
rj885 n16__x_out_2 n18__x_out_2 500e-3
rj886 n15__y_out_0 n16__y_out_0 646.2e-3
rj887 n16__y_out_0 n12__y_out_0 32.21e-3
rj888 n14__y_out_0 n16__y_out_0 500e-3
rj889 n71__i18__net4 n72__i18__net4 500e-3
rj890 n7__ck4 n9__ck4 1.0302
rj891 n12__ck_b n13__ck_b 782.6e-3
rj892 n13__ck_b n6__ck_b 614.6e-3
rj893 n13__ck_b n10__ck_b 588.2e-3
rj894 n463__vddio n464__vddio 333.3e-3
rj895 n465__vddio n466__vddio 333.3e-3
rj896 n467__vddio n468__vddio 333.3e-3
rj897 n12__net11 n11__net11 727.2e-3
rj898 n76__i18__net4 n77__i18__net4 1
rj899 n13__y_out_2 n17__y_out_2 533e-3
rj900 n17__y_out_2 n11__y_out_2 139e-3
rj902 n17__y_out_2 n19__y_out_2 695.3e-3
rj903 n15__x_out_0 n17__x_out_0 533e-3
rj904 n17__x_out_0 n12__x_out_0 143.9e-3
rj906 n17__x_out_0 n19__x_out_0 695.3e-3
rj907 n550__i18__net5 n544__i18__net5 1
rj908 n548__i18__net5 n551__i18__net5 1
rj909 n6__i13__i14__net2 n12__i13__i14__net2 547.5e-3
rj910 n12__i13__i14__net2 n13__i13__i14__net2 174.4e-3
rj911 n12__i13__i14__net2 n4__i13__i14__net2 681.8e-3
rj912 n7__i13__i14__net2 n13__i13__i14__net2 500e-3
rj913 n6__i13__i12__net2 n12__i13__i12__net2 547.5e-3
rj914 n12__i13__i12__net2 n4__i13__i12__net2 681.8e-3
rj915 n12__i13__i12__net2 n10__i13__i12__net2 674.6e-3
rj916 n23__x_out_2 n21__x_out_2 502.5e-3
rj917 n19__y_out_0 n17__y_out_0 502.5e-3
rj918 n78__i18__net4 n79__i18__net4 500e-3
rj919 n16__ck_b n8__ck_b 979.5e-3
rj920 n8__ck_b n14__ck_b 609.3e-3
rj921 n469__vddio n470__vddio 333.3e-3
rj922 n471__vddio n472__vddio 333.3e-3
rj923 n473__vddio n474__vddio 333.3e-3
rj924 n86__i18__net4 n87__i18__net4 500e-3
rj925 n10__ck_buff n9__ck_buff 54.36e-3
rj926 n9__ck_buff n7__ck_buff 1.0137
rj927 n554__i18__net5 n555__i18__net5 1
rj928 n556__i18__net5 n557__i18__net5 1
rj929 n91__i18__net4 n92__i18__net4 1
rj930 n20__i13__a2 n18__i13__a2 321.3e-3
rj931 n18__i13__a2 n12__i13__a2 249.9e-3
rj932 n19__i13__a0 n17__i13__a0 321.3e-3
rj933 n17__i13__a0 n12__i13__a0 249.9e-3
rj934 n6__reset_buff n3__reset_buff 1
rj935 n475__vddio n476__vddio 333.3e-3
rj936 n477__vddio n478__vddio 333.3e-3
rj937 n479__vddio n480__vddio 333.3e-3
rj938 n16__i9__i4__net1 n14__i9__i4__net1 669.1e-3
rj939 n14__i9__i4__net1 n11__i9__i4__net1 1.1446
rj940 n93__i18__net4 n94__i18__net4 1
rj941 n576__i18__net5 n570__i18__net5 1
rj942 n574__i18__net5 n577__i18__net5 1
rj943 n5__i9__i4__net2 n4__i9__i4__net2 1.2876
rj944 n18__x_out_3 n19__x_out_3 642e-3
rj945 n19__x_out_3 n15__x_out_3 524.4e-3
rj946 n17__x_out_3 n19__x_out_3 500e-3
rj947 n17__x_out_1 n18__x_out_1 646.2e-3
rj948 n18__x_out_1 n14__x_out_1 24.35e-3
rj949 n16__x_out_1 n18__x_out_1 500e-3
rj950 n98__i18__net4 n99__i18__net4 500e-3
rj951 n481__vddio n482__vddio 333.3e-3
rj952 n483__vddio n484__vddio 333.3e-3
rj953 n485__vddio n486__vddio 333.3e-3
rj955 n106__i18__net4 n107__i18__net4 500e-3
rj956 n4__reset_b n13__reset_b 488.5e-3
rj957 n13__reset_b n11__reset_b 696.6e-3
rj958 n8__reset_b n13__reset_b 500e-3
rj959 n14__y_out_3 n16__y_out_3 533e-3
rj960 n16__y_out_3 n12__y_out_3 139e-3
rj962 n16__y_out_3 n18__y_out_3 695.3e-3
rj963 n13__y_out_1 n17__y_out_1 533e-3
rj964 n17__y_out_1 n11__y_out_1 143.9e-3
rj966 n17__y_out_1 n19__y_out_1 695.3e-3
rj967 n589__i18__net5 n583__i18__net5 1
rj968 n587__i18__net5 n590__i18__net5 1
rj969 n18__ck_b n17__ck_b 731.9e-3
rj970 n12__ck_buff n11__ck_buff 829e-3
rj971 n6__i13__i15__net2 n12__i13__i15__net2 547.5e-3
rj972 n12__i13__i15__net2 n13__i13__i15__net2 174.4e-3
rj973 n12__i13__i15__net2 n4__i13__i15__net2 681.8e-3
rj974 n7__i13__i15__net2 n13__i13__i15__net2 500e-3
rj975 n6__i13__i13__net2 n12__i13__i13__net2 547.5e-3
rj976 n12__i13__i13__net2 n4__i13__i13__net2 681.8e-3
rj977 n12__i13__i13__net2 n10__i13__i13__net2 674.6e-3
rj978 n22__x_out_3 n20__x_out_3 502.5e-3
rj979 n23__x_out_1 n19__x_out_1 502.5e-3
rj980 n12__net12 n11__net12 727.2e-3
rj981 n108__i18__net4 n109__i18__net4 500e-3
rj982 n487__vddio n488__vddio 333.3e-3
rj983 n489__vddio n490__vddio 333.3e-3
rj984 n491__vddio n492__vddio 333.3e-3
rj985 n116__i18__net4 n117__i18__net4 500e-3
rj986 n593__i18__net5 n594__i18__net5 1
rj987 n595__i18__net5 n596__i18__net5 1
rj988 n118__i18__net4 n119__i18__net4 1
rj989 n17__i13__a3 n16__i13__a3 824.8e-3
rj990 n16__i13__a3 n12__i13__a3 249.9e-3
rj991 n17__i13__a1 n15__i13__a1 824.8e-3
rj992 n15__i13__a1 n12__i13__a1 249.9e-3
rj993 n14__reset_b n6__reset_b 1.7827
rj994 n493__vddio n494__vddio 333.3e-3
rj995 n495__vddio n496__vddio 333.3e-3
rj996 n497__vddio n498__vddio 333.3e-3
rj997 n503__vss n504__vss 166.7e-3
rj998 n505__vss n506__vss 166.7e-3
rj999 n14__i9__i4__net5 n11__i9__i4__net5 1.447
rj1000 n34__ck n35__ck 500e-3
rj1001 n123__i18__net4 n124__i18__net4 500e-3
rj1002 n615__i18__net5 n609__i18__net5 1
rj1003 n613__i18__net5 n616__i18__net5 1
rj1004 n125__i18__net4 n126__i18__net4 500e-3
rj1005 n12__i9__i4__net4 n7__i9__i4__net4 524.3e-3
rj1006 n7__i13__i17__net1 n5__i13__i17__net1 689.4e-3
rj1007 n7__i13__i16__net1 n6__i13__i16__net1 689.4e-3
rj1008 n499__vddio n500__vddio 333.3e-3
rj1009 n501__vddio n502__vddio 333.3e-3
rj1010 n503__vddio n504__vddio 333.3e-3
rj1011 n60__reset n61__reset 250e-3
rj1012 n127__i18__net4 n128__i18__net4 500e-3
rj1013 n13__i9__i4__net4 n9__i9__i4__net4 712.6e-3
rj1014 n622__i18__net5 n628__i18__net5 1
rj1015 n629__i18__net5 n626__i18__net5 1
rj1016 n63__reset n64__reset 250e-3
rj1017 n129__i18__net4 n130__i18__net4 1
rj1018 n505__vddio n506__vddio 333.3e-3
rj1019 n507__vddio n508__vddio 333.3e-3
rj1020 n509__vddio n510__vddio 333.3e-3
rj1021 n15__net13 n11__net13 1.2272
rj1023 n22__ck_buff n14__ck_buff 698.8e-3
rj1024 n25__ck_buff n22__ck_buff 500e-3
rj1025 n132__i18__net4 n131__i18__net4 500e-3
rj1026 n633__i18__net5 n636__i18__net5 500e-3
rj1027 n637__i18__net5 n634__i18__net5 500e-3
rj1028 n25__i13__a2 n26__i13__a2 643.2e-3
rj1029 n26__i13__a2 n23__i13__a2 517.9e-3
rj1030 n23__i13__a2 n22__i13__a2 267.6e-3
rj1031 n24__i13__a2 n26__i13__a2 500e-3
rj1032 n25__i13__a0 n26__i13__a0 643.2e-3
rj1033 n26__i13__a0 n23__i13__a0 517.9e-3
rj1034 n23__i13__a0 n21__i13__a0 267.6e-3
rj1035 n24__i13__a0 n26__i13__a0 500e-3
rj1036 n133__i18__net4 n134__i18__net4 500e-3
rj1037 n511__vddio n512__vddio 333.3e-3
rj1038 n513__vddio n514__vddio 333.3e-3
rj1039 n515__vddio n516__vddio 333.3e-3
rj1040 n10__i9__net1 n11__i9__net1 761.5e-3
rj1041 n8__i9__net1 n11__i9__net1 500e-3
rj1042 n15__net14 n14__net14 727.2e-3
rj1043 n135__i18__net4 n136__i18__net4 500e-3
rj1044 n21__i13__a3 n23__i13__a3 533e-3
rj1045 n23__i13__a3 n19__i13__a3 837.6e-3
rj1046 n19__i13__a3 n18__i13__a3 167.2e-3
rj1047 n23__i13__a3 n24__i13__a3 695.3e-3
rj1048 n21__i13__a1 n23__i13__a1 533e-3
rj1049 n23__i13__a1 n19__i13__a1 837.6e-3
rj1050 n19__i13__a1 n18__i13__a1 167.2e-3
rj1051 n23__i13__a1 n24__i13__a1 695.3e-3
rj1052 n6__i13__i17__i4__net2 n12__i13__i17__i4__net2 547.5e-3
rj1053 n12__i13__i17__i4__net2 n13__i13__i17__i4__net2 190.9e-3
rj1054 n12__i13__i17__i4__net2 n4__i13__i17__i4__net2 700.5e-3
rj1055 n7__i13__i17__i4__net2 n13__i13__i17__i4__net2 500e-3
rj1056 n6__i13__i16__i4__net2 n12__i13__i16__i4__net2 547.5e-3
rj1057 n12__i13__i16__i4__net2 n4__i13__i16__i4__net2 700.5e-3
rj1058 n12__i13__i16__i4__net2 n10__i13__i16__i4__net2 691.1e-3
rj1059 n29__i13__a2 n27__i13__a2 502.5e-3
rj1060 n29__i13__a0 n27__i13__a0 502.5e-3
rj1061 n654__i18__net5 n648__i18__net5 1
rj1062 n652__i18__net5 n655__i18__net5 1
rj1063 n16__ck4 n17__ck4 1
rj1064 n16__reset_buff n17__reset_buff 642.3e-3
rj1065 n17__reset_buff n11__reset_buff 696.6e-3
rj1066 n14__reset_buff n17__reset_buff 500e-3
rj1067 n138__i18__net4 n137__i18__net4 500e-3
rj1068 n517__vddio n518__vddio 333.3e-3
rj1069 n519__vddio n520__vddio 333.3e-3
rj1070 n521__vddio n522__vddio 333.3e-3
rj1071 n5__i9__i1__net1 n4__i9__i1__net1 689.4e-3
rj1072 n4__i9__i1__net1 n2__i9__i1__net1 189.4e-3
rj1073 n139__i18__net4 n140__i18__net4 500e-3
rj1074 n661__i18__net5 n667__i18__net5 1
rj1075 n668__i18__net5 n665__i18__net5 1
rj1076 n16__i13__net1 n11__i13__net1 869.2e-3
rj1077 n17__i13__net12 n16__i13__net12 219.9e-3
rj1078 n16__i13__net12 n12__i13__net12 249.9e-3
rj1079 n19__i13__net2 n17__i13__net2 836.1e-3
rj1080 n17__i13__net2 n14__i13__net2 249.9e-3
rj1081 n13__i13__net11 n9__i13__net11 1.5673
rj1082 n142__i18__net4 n141__i18__net4 500e-3
rj1083 n523__vddio n524__vddio 333.3e-3
rj1084 n525__vddio n526__vddio 333.3e-3
rj1085 n527__vddio n528__vddio 333.3e-3
rj1086 n143__i18__net4 n144__i18__net4 500e-3
rj1087 net4 n2__net4 1
rj1088 net3 n2__net3 1
rj1089 n526__vss n527__vss 1
rj1090 n530__vss n531__vss 1
rj1091 n10__i2__net79 n8__i2__net79 1.3426
rj1092 n10__i1__net79 n8__i1__net79 1.3426
rj1093 n10__i0__net79 n8__i0__net79 1.3426
rj1094 n671__i18__net5 n672__i18__net5 1
rj1095 n673__i18__net5 n674__i18__net5 1
rj1096 n7__i13__i19__net1 n5__i13__i19__net1 689.4e-3
rj1097 n7__i13__i18__net1 n6__i13__i18__net1 689.4e-3
rj1098 n145__i18__net4 n146__i18__net4 500e-3
rj1099 n11__i2__net79 n5__i2__net79 244.8e-3
rj1100 n11__i1__net79 n5__i1__net79 244.8e-3
rj1101 n11__i0__net79 n5__i0__net79 244.8e-3
rj1102 n37__shift n40__shift 749.9e-3
rj1103 n40__shift n41__shift 239.7e-3
rj1104 n41__shift n42__shift 139.1e-3
rj1105 n42__shift n43__shift 201e-3
rj1106 n43__shift n28__shift 211.1e-3
rj1107 n42__shift n44__shift 513.3e-3
rj1108 n44__shift n45__shift 955.7e-3
rj1109 n45__shift n46__shift 239.7e-3
rj1110 n43__shift n30__shift 225.2e-3
rj1111 n28__shift n26__shift 221.7e-3
rj1112 n44__shift n47__shift 86.16e-3
rj1113 n47__shift n48__shift 241.9e-3
rj1114 n46__shift n39__shift 749.9e-3
rj1115 n48__shift n38__shift 752.1e-3
rj1116 n34__shift n40__shift 500e-3
rj1117 n31__shift n41__shift 500e-3
rj1118 n33__shift n45__shift 500e-3
rj1119 n36__shift n46__shift 500e-3
rj1120 n32__shift n47__shift 500e-3
rj1121 n35__shift n48__shift 500e-3
rj1122 n529__vddio n530__vddio 333.3e-3
rj1123 n531__vddio n532__vddio 333.3e-3
rj1124 n533__vddio n534__vddio 333.3e-3
rj1125 n6__r0_buff n4__r0_buff 1
rj1126 n4__r1_buff n6__r1_buff 1
rj1127 n6__r2_buff n4__r2_buff 1
rj1128 n147__i18__net4 n148__i18__net4 500e-3
rj1129 n23__vdd n24__vdd 166.7e-3
rj1130 n693__i18__net5 n687__i18__net5 1
rj1131 n691__i18__net5 n694__i18__net5 1
rj1132 n149__i18__net4 n150__i18__net4 125e-3
rj1134 n606__vss n608__vss 944.2e-3
rj1136 n608__vss n610__vss 1.0491
rj1138 n610__vss n612__vss 1.0491
rj1139 n612__vss n613__vss 25e-3
rj1140 n545__vss n606__vss 31.25e-3
rj1141 n562__vss n608__vss 25e-3
rj1142 n581__vss n610__vss 25e-3
rj1143 n598__vss n612__vss 25e-3
rj1145 n626__vddio n628__vddio 944.2e-3
rj1147 n628__vddio n630__vddio 1.0491
rj1149 n630__vddio n632__vddio 1.0491
rj1150 n632__vddio n558__vddio 25e-3
rj1151 n543__vddio n626__vddio 31.25e-3
rj1152 n548__vddio n628__vddio 25e-3
rj1153 n553__vddio n630__vddio 25e-3
rj1154 n614__vss n536__vss 333.3e-3
rj1155 n537__vddio n633__vddio 333.3e-3
rj1156 n634__vddio n539__vddio 333.3e-3
rj1157 n541__vddio n635__vddio 333.3e-3
rj1158 n19__i13__net1 n20__i13__net1 643.2e-3
rj1159 n20__i13__net1 n17__i13__net1 517.9e-3
rj1160 n17__i13__net1 n15__i13__net1 369.9e-3
rj1161 n18__i13__net1 n20__i13__net1 500e-3
rj1162 n23__i13__net2 n24__i13__net2 643.2e-3
rj1163 n24__i13__net2 n21__i13__net2 517.9e-3
rj1164 n21__i13__net2 n20__i13__net2 267.6e-3
rj1165 n22__i13__net2 n24__i13__net2 500e-3
rj1166 n17__i13__net11 n19__i13__net11 533e-3
rj1167 n19__i13__net11 n15__i13__net11 837.6e-3
rj1168 n15__i13__net11 n14__i13__net11 167.2e-3
rj1169 n19__i13__net11 n20__i13__net11 695.3e-3
rj1170 n21__i13__net12 n23__i13__net12 533e-3
rj1171 n23__i13__net12 n19__i13__net12 837.6e-3
rj1172 n19__i13__net12 n18__i13__net12 281e-3
rj1173 n23__i13__net12 n24__i13__net12 695.3e-3
rj1174 n6__i13__i19__i4__net2 n12__i13__i19__i4__net2 547.5e-3
rj1175 n12__i13__i19__i4__net2 n13__i13__i19__i4__net2 190.9e-3
rj1176 n12__i13__i19__i4__net2 n4__i13__i19__i4__net2 700.5e-3
rj1177 n7__i13__i19__i4__net2 n13__i13__i19__i4__net2 500e-3
rj1178 n6__i13__i18__i4__net2 n12__i13__i18__i4__net2 547.5e-3
rj1179 n12__i13__i18__i4__net2 n4__i13__i18__i4__net2 700.5e-3
rj1180 n12__i13__i18__i4__net2 n10__i13__i18__i4__net2 691.1e-3
rj1181 n23__i13__net1 n21__i13__net1 502.5e-3
rj1182 n27__i13__net2 n25__i13__net2 502.5e-3
rj1183 n31__i18__net3 n32__i18__net3 500e-3
rj1184 n154__i18__net4 n159__i18__net4 1
rj1185 n160__i18__net4 n157__i18__net4 1
rj1186 n34__i18__net3 n33__i18__net3 500e-3
rj1187 n19__i13__net18 n18__i13__net18 724.7e-3
rj1188 n18__i13__net18 n14__i13__net18 249.9e-3
rj1189 n9__r0 n7__r0 628e-3
rj1190 n7__r0 n4__r0 249.9e-3
rj1191 n13__i13__net7 n9__i13__net7 1.5698
rj1192 n37__i18__net3 n35__i18__net3 500e-3
rj1193 n10__i13__net17 n5__i13__net17 1.664
rj1194 n38__ck_b n35__ck_b 975.5e-3
rj1195 n35__ck_b n32__ck_b 1.231
rj1196 n39__ck_b n36__ck_b 975.5e-3
rj1197 n36__ck_b n33__ck_b 1.231
rj1198 n40__ck_b n37__ck_b 975.5e-3
rj1199 n37__ck_b n34__ck_b 731e-3
rj1200 n170__i18__net4 n165__i18__net4 1
rj1201 n168__i18__net4 n171__i18__net4 1
rj1202 n41__ck_buff n38__ck_buff 575.6e-3
rj1203 n38__ck_buff n36__ck_buff 971.1e-3
rj1204 n44__ck_buff n39__ck_buff 575.6e-3
rj1205 n39__ck_buff n34__ck_buff 968.7e-3
rj1206 n45__ck_buff n40__ck_buff 575.6e-3
rj1207 n40__ck_buff n35__ck_buff 471.1e-3
rj1208 n36__i18__net3 n38__i18__net3 500e-3
rj1209 n9__i13__net17 n11__i13__net17 570.1e-3
rj1210 n7__i13__i20__net1 n5__i13__i20__net1 689.4e-3
rj1211 n6__i13__net3 n5__i13__net3 689.4e-3
rj1212 n39__i18__net3 n40__i18__net3 1
rj1213 n30__reset_buff n26__reset_buff 2.0576
rj1214 n31__reset_buff n27__reset_buff 2.5576
rj1215 n32__reset_buff n29__reset_buff 2.0576
rj1216 n175__i18__net4 n178__i18__net4 500e-3
rj1217 n179__i18__net4 n176__i18__net4 500e-3
rj1218 n16__i2__net74 n15__i2__net74 711.4e-3
rj1219 n15__i2__net74 n11__i2__net74 1.1023
rj1220 n16__i1__net74 n15__i1__net74 711.4e-3
rj1221 n15__i1__net74 n11__i1__net74 1.1023
rj1222 n16__i0__net74 n15__i0__net74 711.4e-3
rj1223 n15__i0__net74 n11__i0__net74 1.1023
rj1224 n10__i13__net23 n5__i13__net23 841.8e-3
rj1225 n41__i18__net3 n42__i18__net3 500e-3
rj1226 n4__r2 n2__r2 1.0974
rj1227 n5__i2__net75 n4__i2__net75 1.2876
rj1228 n5__i1__net75 n4__i1__net75 1.2876
rj1229 n5__i0__net75 n4__i0__net75 1.2876
rj1230 n43__i18__net3 n44__i18__net3 500e-3
rj1231 n192__i18__net4 n187__i18__net4 1
rj1232 n190__i18__net4 n193__i18__net4 1
rj1233 n24__i13__net18 n25__i13__net18 143.2e-3
rj1234 n25__i13__net18 n20__i13__net18 517.9e-3
rj1235 n20__i13__net18 n21__i13__net18 365.1e-3
rj1236 n22__i13__net18 n25__i13__net18 500e-3
rj1237 n45__i18__net3 n47__i18__net3 500e-3
rj1238 n44__ck_b n41__ck_b 731.9e-3
rj1239 n45__ck_b n42__ck_b 731.9e-3
rj1240 n46__ck_b n43__ck_b 731.9e-3
rj1241 n47__ck_buff n42__ck_buff 829e-3
rj1242 n48__ck_buff n43__ck_buff 829e-3
rj1243 n49__ck_buff n46__ck_buff 829e-3
rj1244 n48__i18__net3 n46__i18__net3 500e-3
rj1245 n17__i13__net7 n19__i13__net7 533e-3
rj1246 n19__i13__net7 n14__i13__net7 837.6e-3
rj1247 n14__i13__net7 n15__i13__net7 167.2e-3
rj1248 n19__i13__net7 n20__i13__net7 695.3e-3
rj1249 n203__i18__net4 n198__i18__net4 1
rj1250 n201__i18__net4 n204__i18__net4 1
rj1251 n6__i13__i20__i4__net2 n12__i13__i20__i4__net2 547.5e-3
rj1252 n12__i13__i20__i4__net2 n13__i13__i20__i4__net2 190.9e-3
rj1253 n12__i13__i20__i4__net2 n4__i13__i20__i4__net2 700.5e-3
rj1254 n7__i13__i20__i4__net2 n13__i13__i20__i4__net2 500e-3
rj1255 n27__i13__net18 n23__i13__net18 502.5e-3
rj1256 n49__i18__net3 n50__i18__net3 1
rj1258 n1298__vss n1300__vss 681.9e-3
rj1259 n1300__vss n1301__vss 25e-3
rj1260 n625__vss n1298__vss 83.33e-3
rj1261 n628__vss n1300__vss 25e-3
rj1263 n964__vddio n966__vddio 681.9e-3
rj1264 n966__vddio n642__vddio 25e-3
rj1265 n639__vddio n964__vddio 83.33e-3
rj1266 n25__reset_b n22__reset_b 3.2894
rj1267 n26__reset_b n23__reset_b 3.2894
rj1268 n27__reset_b n24__reset_b 2.7894
rj1269 n14__i2__net76 n11__i2__net76 1.447
rj1270 n14__i1__net76 n11__i1__net76 1.447
rj1271 n14__i0__net76 n11__i0__net76 1.447
rj1272 n6__i13__net23 n11__i13__net23 2.416e-3
rj1273 n12__r1 n8__r1 240.5e-3
rj1275 n12__i2__net77 n7__i2__net77 524.3e-3
rj1276 n12__i1__net77 n7__i1__net77 524.3e-3
rj1277 n12__i0__net77 n7__i0__net77 524.3e-3
rj1278 n13__i2__net77 n9__i2__net77 712.6e-3
rj1279 n13__i1__net77 n9__i1__net77 712.6e-3
rj1280 n13__i0__net77 n9__i0__net77 712.6e-3
rj1281 n8__i12__bio n4__i12__bio 910e-3
rj1285 n25__serial_out n22__serial_out 1.2102
rj1286 n16__net4 n13__net4 1.2102
rj1287 n14__net3 n12__net3 1.2102
rj1288 n1302__vss n710__vss 90.91e-3
rj1289 n661__vddio n967__vddio 90.91e-3
rj1290 n5__i12__bcore_bar n16__i12__bcore_bar 682e-3
rj1291 n16__i12__bcore_bar i12__bcore_bar 687.9e-3
rj1292 n3__i12__bcore_bar n16__i12__bcore_bar 500e-3
rj1293 n12__serial_out_b_high n11__serial_out_b_high 380.8e-3
rj1294 n11__serial_out_b_high n14__serial_out_b_high 2.196e-3
rj1295 n11__serial_out_b_high n7__serial_out_b_high 593.1e-3
rj1296 n15__r1 n13__r1 500e-3
rj1297 n14__r0 n15__r0 500e-3
rj1298 n10__r2 n9__r2 500e-3
rj1299 n1303__vss n1003__vss 166.7e-3
rj1300 n680__vddio n968__vddio 166.7e-3
rj1301 n31__vdd n419__vdd 83.33e-3
rj1302 n420__vdd n131__vdd 166.7e-3
rj1303 n24__serial_out n26__serial_out 391.1e-3
rj1304 n26__serial_out n27__serial_out 1.1573
rj1305 n27__serial_out n28__serial_out 160.4e-3
rj1306 n28__serial_out n1__serial_out 660.4e-3
rj1307 n5__serial_out n27__serial_out 500e-3
rj1308 n3__serial_out n28__serial_out 500e-3
rj1309 n15__serial_out_b_high n13__serial_out_b_high 500e-3
rj1310 n684__vddio n969__vddio 166.7e-3
rj1311 n970__vddio n670__vddio 83.33e-3
rj1316 n688__vddio n975__vddio 166.7e-3
rj1317 n12__r0_buff n15__r0_buff 1
rj1318 n16__r2_buff n10__r2_buff 1
rj1319 n12__r1_buff n15__r1_buff 1
rj1320 n1016__vss n1304__vss 83.33e-3
rj1325 n8__serial_out_b_high_buff n4__serial_out_b_high_buff 2.7978
rk1 n2__i18__net5 n46__i18__net5 45
rk2 n7__r_out n8__r_out 8.6557
rk3 n8__r_out n9__r_out 1.541
rk4 n9__r_out n1__r_out 40.59e-3
rk6 n7__r_out n8__r_out 3.75
rk7 n7__r_out n9__r_out 3.75
rk8 n11__r_out n12__r_out 8.8496
rk9 n12__r_out n4__r_out 119.8e-3
rk10 n4__r_out n13__r_out 1.4232
rk11 n13__r_out n11__r_out 4.641
rk12 n11__r_out n12__r_out 3.1
rk13 n11__r_out n13__r_out 3.1
rk14 n5__i18__net5 n48__i18__net5 45.5
rk15 n8__i18__net5 n56__i18__net5 45
rk16 n14__r_out n15__r_out 8.6557
rk17 n15__r_out n16__r_out 1.541
rk18 n16__r_out n17__r_out 28.99e-3
rk20 n14__r_out n15__r_out 3.75
rk21 n14__r_out n16__r_out 3.75
rk22 n19__r_out n20__r_out 8.8496
rk23 n20__r_out n21__r_out 105.1e-3
rk24 n21__r_out n22__r_out 1.4342
rk25 n22__r_out n19__r_out 4.641
rk26 n19__r_out n20__r_out 3.1
rk27 n19__r_out n22__r_out 3.1
rk28 n11__i18__net5 n58__i18__net5 45.5
rk29 n14__i18__net5 n66__i18__net5 45
rk30 n31__r_out n32__r_out 8.6557
rk31 n32__r_out n33__r_out 1.541
rk32 n33__r_out n27__r_out 37.69e-3
rk34 n31__r_out n32__r_out 3.75
rk35 n31__r_out n33__r_out 3.75
rk36 n35__r_out n36__r_out 8.8496
rk37 n36__r_out n30__r_out 114.7e-3
rk38 n30__r_out n37__r_out 1.4246
rk39 n37__r_out n35__r_out 4.641
rk40 n35__r_out n36__r_out 3.1
rk41 n35__r_out n37__r_out 3.1
rk42 n17__i18__net5 n71__i18__net5 45.5
rk43 n20__i18__net5 n76__i18__net5 45
rk44 n46__r_out n47__r_out 8.6557
rk45 n47__r_out n48__r_out 1.541
rk46 n48__r_out n40__r_out 40.59e-3
rk48 n46__r_out n47__r_out 3.75
rk49 n46__r_out n48__r_out 3.75
rk50 n50__r_out n51__r_out 8.8496
rk51 n51__r_out n43__r_out 119.8e-3
rk52 n43__r_out n52__r_out 1.4232
rk53 n52__r_out n50__r_out 4.641
rk54 n50__r_out n51__r_out 3.1
rk55 n50__r_out n52__r_out 3.1
rk56 n23__i18__net5 n81__i18__net5 45.5
rk57 n26__i18__net5 n83__i18__net5 45.5
rk58 n57__r_out n58__r_out 8.6557
rk59 n58__r_out n59__r_out 1.541
rk60 n59__r_out n53__r_out 28.99e-3
rk62 n57__r_out n58__r_out 3.75
rk63 n57__r_out n59__r_out 3.75
rk64 n61__r_out n62__r_out 8.8496
rk65 n62__r_out n56__r_out 105.1e-3
rk66 n56__r_out n63__r_out 1.4342
rk67 n63__r_out n61__r_out 4.641
rk68 n61__r_out n62__r_out 3.1
rk69 n61__r_out n63__r_out 3.1
rk70 n29__i18__net5 n88__i18__net5 45.5
rk71 n32__i18__net5 n93__i18__net5 45
rk72 n72__r_out n73__r_out 8.6557
rk73 n73__r_out n74__r_out 1.541
rk74 n74__r_out n66__r_out 40.59e-3
rk76 n72__r_out n73__r_out 3.75
rk77 n72__r_out n74__r_out 3.75
rk78 n76__r_out n77__r_out 8.8496
rk79 n77__r_out n69__r_out 119.8e-3
rk80 n69__r_out n78__r_out 1.4232
rk81 n78__r_out n76__r_out 4.641
rk82 n76__r_out n77__r_out 3.1
rk83 n76__r_out n78__r_out 3.1
rk84 n35__i18__net5 n98__i18__net5 45.5
rk85 n38__i18__net5 n106__i18__net5 45
rk86 n79__r_out n80__r_out 8.6557
rk87 n80__r_out n81__r_out 1.541
rk88 n81__r_out n82__r_out 28.99e-3
rk90 n79__r_out n80__r_out 3.75
rk91 n79__r_out n81__r_out 3.75
rk92 n84__r_out n85__r_out 8.8496
rk93 n85__r_out n86__r_out 107e-3
rk94 n86__r_out n87__r_out 1.4361
rk95 n87__r_out n84__r_out 4.641
rk96 n84__r_out n85__r_out 3.1
rk97 n84__r_out n87__r_out 3.1
rk98 n41__i18__net5 n109__i18__net5 45
rk99 n44__i18__net5 n113__i18__net5 45
rk100 n98__r_out n99__r_out 8.6557
rk101 n99__r_out n100__r_out 1.541
rk102 n100__r_out n92__r_out 37.69e-3
rk104 n98__r_out n99__r_out 3.75
rk105 n98__r_out n100__r_out 3.75
rk106 n102__r_out n103__r_out 8.8496
rk107 n103__r_out n95__r_out 116.6e-3
rk108 n95__r_out n104__r_out 1.4265
rk109 n104__r_out n102__r_out 4.641
rk110 n102__r_out n103__r_out 3.1
rk111 n102__r_out n104__r_out 3.1
rk112 n51__i18__net5 n119__i18__net5 45
rk113 n54__i18__net5 n126__i18__net5 45
rk114 n111__r_out n112__r_out 8.6557
rk115 n112__r_out n113__r_out 1.541
rk116 n113__r_out n105__r_out 40.59e-3
rk118 n111__r_out n112__r_out 3.75
rk119 n111__r_out n113__r_out 3.75
rk120 n115__r_out n116__r_out 8.8496
rk121 n116__r_out n108__r_out 119.8e-3
rk122 n108__r_out n117__r_out 1.4232
rk123 n117__r_out n115__r_out 4.641
rk124 n115__r_out n116__r_out 3.1
rk125 n115__r_out n117__r_out 3.1
rk126 n61__i18__net5 n128__i18__net5 45.5
rk127 n64__i18__net5 n133__i18__net5 45
rk128 n124__r_out n125__r_out 8.6557
rk129 n125__r_out n126__r_out 1.541
rk130 n126__r_out n118__r_out 28.99e-3
rk132 n124__r_out n125__r_out 3.75
rk133 n124__r_out n126__r_out 3.75
rk134 n128__r_out n129__r_out 8.8496
rk135 n129__r_out n121__r_out 107e-3
rk136 n121__r_out n130__r_out 1.4361
rk137 n130__r_out n128__r_out 4.641
rk138 n128__r_out n129__r_out 3.1
rk139 n128__r_out n130__r_out 3.1
rk140 n69__i18__net5 n141__i18__net5 45.5
rk141 n74__i18__net5 n146__i18__net5 45.5
rk142 n131__r_out n132__r_out 8.6557
rk143 n132__r_out n133__r_out 1.541
rk144 n133__r_out n134__r_out 40.59e-3
rk146 n131__r_out n132__r_out 3.75
rk147 n131__r_out n133__r_out 3.75
rk148 n136__r_out n137__r_out 8.8496
rk149 n137__r_out n138__r_out 119.8e-3
rk150 n138__r_out n139__r_out 1.4232
rk151 n139__r_out n136__r_out 4.641
rk152 n136__r_out n137__r_out 3.1
rk153 n136__r_out n139__r_out 3.1
rk154 n79__i18__net5 n151__i18__net5 45.5
rk155 n86__i18__net5 n156__i18__net5 45
rk156 n144__r_out n145__r_out 8.6557
rk157 n145__r_out n146__r_out 1.541
rk158 n146__r_out n147__r_out 28.99e-3
rk160 n144__r_out n145__r_out 3.75
rk161 n144__r_out n146__r_out 3.75
rk162 n149__r_out n150__r_out 8.8496
rk163 n150__r_out n151__r_out 105.1e-3
rk164 n151__r_out n152__r_out 1.4342
rk165 n152__r_out n149__r_out 4.641
rk166 n149__r_out n150__r_out 3.1
rk167 n149__r_out n152__r_out 3.1
rk168 n91__i18__net5 n158__i18__net5 45.5
rk169 n96__i18__net5 n163__i18__net5 45.5
rk170 n161__r_out n162__r_out 8.6557
rk171 n162__r_out n163__r_out 1.541
rk172 n163__r_out n157__r_out 37.69e-3
rk174 n161__r_out n162__r_out 3.75
rk175 n161__r_out n163__r_out 3.75
rk176 n165__r_out n166__r_out 8.8496
rk177 n166__r_out n160__r_out 114.7e-3
rk178 n160__r_out n167__r_out 1.4246
rk179 n167__r_out n165__r_out 4.641
rk180 n165__r_out n166__r_out 3.1
rk181 n165__r_out n167__r_out 3.1
rk182 n101__i18__net5 n168__i18__net5 45.5
rk183 n104__i18__net5 n176__i18__net5 45
rk184 n176__r_out n177__r_out 8.6557
rk185 n177__r_out n178__r_out 1.541
rk186 n178__r_out n170__r_out 40.59e-3
rk188 n176__r_out n177__r_out 3.75
rk189 n176__r_out n178__r_out 3.75
rk190 n180__r_out n181__r_out 8.8496
rk191 n181__r_out n173__r_out 119.8e-3
rk192 n173__r_out n182__r_out 1.4232
rk193 n182__r_out n180__r_out 4.641
rk194 n180__r_out n181__r_out 3.1
rk195 n180__r_out n182__r_out 3.1
rk196 n111__i18__net5 n178__i18__net5 45.5
rk197 n116__i18__net5 n183__i18__net5 45
rk198 n187__r_out n188__r_out 8.6557
rk199 n188__r_out n189__r_out 1.541
rk200 n189__r_out n183__r_out 28.99e-3
rk202 n187__r_out n188__r_out 3.75
rk203 n187__r_out n189__r_out 3.75
rk204 n191__r_out n192__r_out 8.8496
rk205 n192__r_out n186__r_out 105.1e-3
rk206 n186__r_out n193__r_out 1.4342
rk207 n193__r_out n191__r_out 4.641
rk208 n191__r_out n192__r_out 3.1
rk209 n191__r_out n193__r_out 3.1
rk210 n121__i18__net5 n191__i18__net5 45.5
rk211 n124__i18__net5 n196__i18__net5 45
rk212 n202__r_out n203__r_out 8.6557
rk213 n203__r_out n204__r_out 1.541
rk214 n204__r_out n196__r_out 40.59e-3
rk216 n202__r_out n203__r_out 3.75
rk217 n202__r_out n204__r_out 3.75
rk218 n206__r_out n207__r_out 8.8496
rk219 n207__r_out n199__r_out 119.8e-3
rk220 n199__r_out n208__r_out 1.4232
rk221 n208__r_out n206__r_out 4.641
rk222 n206__r_out n207__r_out 3.1
rk223 n206__r_out n208__r_out 3.1
rk224 n130__i18__net5 n198__i18__net5 45.5
rk225 n136__i18__net5 n206__i18__net5 45
rk226 n209__r_out n210__r_out 8.6557
rk227 n210__r_out n211__r_out 1.541
rk228 n211__r_out n212__r_out 28.99e-3
rk230 n209__r_out n210__r_out 3.75
rk231 n209__r_out n211__r_out 3.75
rk232 n214__r_out n215__r_out 8.8496
rk233 n215__r_out n216__r_out 107e-3
rk234 n216__r_out n217__r_out 1.4361
rk235 n217__r_out n214__r_out 4.641
rk236 n214__r_out n215__r_out 3.1
rk237 n214__r_out n217__r_out 3.1
rk238 n139__i18__net5 n211__i18__net5 45.5
rk239 n144__i18__net5 n213__i18__net5 45.5
rk240 n228__r_out n229__r_out 8.6557
rk241 n229__r_out n230__r_out 1.541
rk242 n230__r_out n222__r_out 37.69e-3
rk244 n228__r_out n229__r_out 3.75
rk245 n228__r_out n230__r_out 3.75
rk246 n232__r_out n233__r_out 8.8496
rk247 n233__r_out n225__r_out 116.6e-3
rk248 n225__r_out n234__r_out 1.4265
rk249 n234__r_out n232__r_out 4.641
rk250 n232__r_out n233__r_out 3.1
rk251 n232__r_out n234__r_out 3.1
rk252 n149__i18__net5 n221__i18__net5 45.5
rk253 n154__i18__net5 n226__i18__net5 45
rk254 n241__r_out n242__r_out 8.6557
rk255 n242__r_out n243__r_out 1.541
rk256 n243__r_out n235__r_out 40.59e-3
rk258 n241__r_out n242__r_out 3.75
rk259 n241__r_out n243__r_out 3.75
rk260 n245__r_out n246__r_out 8.8496
rk261 n246__r_out n238__r_out 119.8e-3
rk262 n238__r_out n247__r_out 1.4232
rk263 n247__r_out n245__r_out 4.641
rk264 n245__r_out n246__r_out 3.1
rk265 n245__r_out n247__r_out 3.1
rk266 n161__i18__net5 n231__i18__net5 45.5
rk267 n165__i18__net5 n233__i18__net5 45.5
rk268 n254__r_out n255__r_out 8.6557
rk269 n255__r_out n256__r_out 1.541
rk270 n256__r_out n248__r_out 28.99e-3
rk272 n254__r_out n255__r_out 3.75
rk273 n254__r_out n256__r_out 3.75
rk274 n258__r_out n259__r_out 8.8496
rk275 n259__r_out n251__r_out 107e-3
rk276 n251__r_out n260__r_out 1.4361
rk277 n260__r_out n258__r_out 4.641
rk278 n258__r_out n259__r_out 3.1
rk279 n258__r_out n260__r_out 3.1
rk280 n171__i18__net5 n238__i18__net5 45.5
rk281 n174__i18__net5 n243__i18__net5 45
rk282 n267__r_out n268__r_out 8.6557
rk283 n268__r_out n269__r_out 1.541
rk284 n269__r_out n261__r_out 40.59e-3
rk286 n267__r_out n268__r_out 3.75
rk287 n267__r_out n269__r_out 3.75
rk288 n271__r_out n272__r_out 8.8496
rk289 n272__r_out n264__r_out 119.8e-3
rk290 n264__r_out n273__r_out 1.4232
rk291 n273__r_out n271__r_out 4.641
rk292 n271__r_out n272__r_out 3.1
rk293 n271__r_out n273__r_out 3.1
rk294 n180__i18__net5 n248__i18__net5 45.5
rk295 n186__i18__net5 n256__i18__net5 45
rk296 n274__r_out n275__r_out 8.6557
rk297 n275__r_out n276__r_out 1.541
rk298 n276__r_out n277__r_out 28.99e-3
rk300 n274__r_out n275__r_out 3.75
rk301 n274__r_out n276__r_out 3.75
rk302 n279__r_out n280__r_out 8.8496
rk303 n280__r_out n281__r_out 107e-3
rk304 n281__r_out n282__r_out 1.4361
rk305 n282__r_out n279__r_out 4.641
rk306 n279__r_out n280__r_out 3.1
rk307 n279__r_out n282__r_out 3.1
rk308 n189__i18__net5 n261__i18__net5 45.5
rk309 n194__i18__net5 n263__i18__net5 45
rk310 n293__r_out n294__r_out 8.6557
rk311 n294__r_out n295__r_out 1.541
rk312 n295__r_out n287__r_out 37.69e-3
rk314 n293__r_out n294__r_out 3.75
rk315 n293__r_out n295__r_out 3.75
rk316 n297__r_out n298__r_out 8.8496
rk317 n298__r_out n290__r_out 116.6e-3
rk318 n290__r_out n299__r_out 1.4265
rk319 n299__r_out n297__r_out 4.641
rk320 n297__r_out n298__r_out 3.1
rk321 n297__r_out n299__r_out 3.1
rk322 n200__i18__net5 n271__i18__net5 45.5
rk323 n204__i18__net5 n273__i18__net5 45
rk324 n306__r_out n307__r_out 8.6557
rk325 n307__r_out n308__r_out 1.541
rk326 n308__r_out n300__r_out 40.59e-3
rk328 n306__r_out n307__r_out 3.75
rk329 n306__r_out n308__r_out 3.75
rk330 n310__r_out n311__r_out 8.8496
rk331 n311__r_out n303__r_out 119.8e-3
rk332 n303__r_out n312__r_out 1.4232
rk333 n312__r_out n310__r_out 4.641
rk334 n310__r_out n311__r_out 3.1
rk335 n310__r_out n312__r_out 3.1
rk336 n209__i18__net5 n281__i18__net5 45.5
rk337 n215__i18__net5 n286__i18__net5 45
rk338 n319__r_out n320__r_out 8.6557
rk339 n320__r_out n321__r_out 1.541
rk340 n321__r_out n313__r_out 28.99e-3
rk342 n319__r_out n320__r_out 3.75
rk343 n319__r_out n321__r_out 3.75
rk344 n323__r_out n324__r_out 8.8496
rk345 n324__r_out n316__r_out 107e-3
rk346 n316__r_out n325__r_out 1.4361
rk347 n325__r_out n323__r_out 4.641
rk348 n323__r_out n324__r_out 3.1
rk349 n323__r_out n325__r_out 3.1
rk350 n219__i18__net5 n291__i18__net5 45.5
rk351 n224__i18__net5 n296__i18__net5 45
rk352 n332__r_out n333__r_out 8.6557
rk353 n333__r_out n334__r_out 1.541
rk354 n334__r_out n326__r_out 40.59e-3
rk356 n332__r_out n333__r_out 3.75
rk357 n332__r_out n334__r_out 3.75
rk358 n336__r_out n337__r_out 8.8496
rk359 n337__r_out n329__r_out 119.8e-3
rk360 n329__r_out n338__r_out 1.4232
rk361 n338__r_out n336__r_out 4.641
rk362 n336__r_out n337__r_out 3.1
rk363 n336__r_out n338__r_out 3.1
rk364 n229__i18__net5 n301__i18__net5 45.5
rk365 n236__i18__net5 n306__i18__net5 45
rk366 n339__r_out n340__r_out 8.6557
rk367 n340__r_out n341__r_out 1.541
rk368 n341__r_out n342__r_out 28.99e-3
rk370 n339__r_out n340__r_out 3.75
rk371 n339__r_out n341__r_out 3.75
rk372 n344__r_out n345__r_out 8.8496
rk373 n345__r_out n346__r_out 105.1e-3
rk374 n346__r_out n347__r_out 1.4342
rk375 n347__r_out n344__r_out 4.641
rk376 n344__r_out n345__r_out 3.1
rk377 n344__r_out n347__r_out 3.1
rk378 n241__i18__net5 n308__i18__net5 45.5
rk379 n246__i18__net5 n316__i18__net5 45
rk380 n356__r_out n357__r_out 8.6557
rk381 n357__r_out n358__r_out 1.541
rk382 n358__r_out n352__r_out 37.69e-3
rk384 n356__r_out n357__r_out 3.75
rk385 n356__r_out n358__r_out 3.75
rk386 n360__r_out n361__r_out 8.8496
rk387 n361__r_out n355__r_out 114.7e-3
rk388 n355__r_out n362__r_out 1.4246
rk389 n362__r_out n360__r_out 4.641
rk390 n360__r_out n361__r_out 3.1
rk391 n360__r_out n362__r_out 3.1
rk392 n251__i18__net5 n318__i18__net5 45.5
rk393 n254__i18__net5 n323__i18__net5 45
rk394 n371__r_out n372__r_out 8.6557
rk395 n372__r_out n373__r_out 1.541
rk396 n373__r_out n365__r_out 40.59e-3
rk398 n371__r_out n372__r_out 3.75
rk399 n371__r_out n373__r_out 3.75
rk400 n375__r_out n376__r_out 8.8496
rk401 n376__r_out n368__r_out 119.8e-3
rk402 n368__r_out n377__r_out 1.4232
rk403 n377__r_out n375__r_out 4.641
rk404 n375__r_out n376__r_out 3.1
rk405 n375__r_out n377__r_out 3.1
rk406 n259__i18__net5 n331__i18__net5 45.5
rk407 n266__i18__net5 n333__i18__net5 45
rk408 n382__r_out n383__r_out 8.6557
rk409 n383__r_out n384__r_out 1.541
rk410 n384__r_out n378__r_out 28.99e-3
rk412 n382__r_out n383__r_out 3.75
rk413 n382__r_out n384__r_out 3.75
rk414 n386__r_out n387__r_out 8.8496
rk415 n387__r_out n381__r_out 105.1e-3
rk416 n381__r_out n388__r_out 1.4342
rk417 n388__r_out n386__r_out 4.641
rk418 n386__r_out n387__r_out 3.1
rk419 n386__r_out n388__r_out 3.1
rk420 n269__i18__net5 n341__i18__net5 45.5
rk421 n276__i18__net5 n343__i18__net5 45
rk422 n395__r_out n396__r_out 8.6557
rk423 n396__r_out n397__r_out 1.541
rk424 n397__r_out n391__r_out 40.59e-3
rk426 n395__r_out n396__r_out 3.75
rk427 n395__r_out n397__r_out 3.75
rk428 n399__r_out n400__r_out 8.8496
rk429 n400__r_out n394__r_out 119.8e-3
rk430 n394__r_out n401__r_out 1.4232
rk431 n401__r_out n399__r_out 4.641
rk432 n399__r_out n400__r_out 3.1
rk433 n399__r_out n401__r_out 3.1
rk434 n279__i18__net5 n351__i18__net5 45.5
rk435 n284__i18__net5 n353__i18__net5 45
rk436 n404__r_out n405__r_out 8.6557
rk437 n405__r_out n406__r_out 1.541
rk438 n406__r_out n407__r_out 28.99e-3
rk440 n404__r_out n405__r_out 3.75
rk441 n404__r_out n406__r_out 3.75
rk442 n409__r_out n410__r_out 8.8496
rk443 n410__r_out n411__r_out 107e-3
rk444 n411__r_out n412__r_out 1.4361
rk445 n412__r_out n409__r_out 4.641
rk446 n409__r_out n410__r_out 3.1
rk447 n409__r_out n412__r_out 3.1
rk448 n289__i18__net5 n358__i18__net5 45.5
rk449 n294__i18__net5 n363__i18__net5 45
rk450 n417__r_out n418__r_out 8.6557
rk451 n418__r_out n419__r_out 1.541
rk452 n419__r_out n420__r_out 37.69e-3
rk454 n417__r_out n418__r_out 3.75
rk455 n417__r_out n419__r_out 3.75
rk456 n422__r_out n423__r_out 8.8496
rk457 n423__r_out n424__r_out 116.6e-3
rk458 n424__r_out n425__r_out 1.4265
rk459 n425__r_out n422__r_out 4.641
rk460 n422__r_out n423__r_out 3.1
rk461 n422__r_out n425__r_out 3.1
rk462 n299__i18__net5 n371__i18__net5 45.5
rk463 n304__i18__net5 n373__i18__net5 45.5
rk464 n438__r_out n439__r_out 8.6557
rk465 n439__r_out n440__r_out 1.541
rk466 n440__r_out n432__r_out 40.59e-3
rk468 n438__r_out n439__r_out 3.75
rk469 n438__r_out n440__r_out 3.75
rk470 n442__r_out n443__r_out 8.8496
rk471 n443__r_out n435__r_out 119.8e-3
rk472 n435__r_out n444__r_out 1.4232
rk473 n444__r_out n442__r_out 4.641
rk474 n442__r_out n443__r_out 3.1
rk475 n442__r_out n444__r_out 3.1
rk476 n311__i18__net5 n381__i18__net5 45.5
rk477 n314__i18__net5 n383__i18__net5 45.5
rk478 n445__r_out n446__r_out 8.6557
rk479 n446__r_out n447__r_out 1.541
rk480 n447__r_out n448__r_out 28.99e-3
rk482 n445__r_out n446__r_out 3.75
rk483 n445__r_out n447__r_out 3.75
rk484 n450__r_out n451__r_out 8.8496
rk485 n451__r_out n452__r_out 107e-3
rk486 n452__r_out n453__r_out 1.4361
rk487 n453__r_out n450__r_out 4.641
rk488 n450__r_out n451__r_out 3.1
rk489 n450__r_out n453__r_out 3.1
rk490 n321__i18__net5 n388__i18__net5 45.5
rk491 n326__i18__net5 n393__i18__net5 45.5
rk492 n461__r_out n462__r_out 8.6557
rk493 n462__r_out n463__r_out 1.541
rk494 n463__r_out n464__r_out 43.48e-3
rk496 n461__r_out n462__r_out 3.75
rk497 n461__r_out n463__r_out 3.75
rk498 n466__r_out n467__r_out 8.8496
rk499 n467__r_out n468__r_out 119.8e-3
rk500 n468__r_out n469__r_out 1.4232
rk501 n469__r_out n466__r_out 4.641
rk502 n466__r_out n467__r_out 3.1
rk503 n466__r_out n469__r_out 3.1
rk504 n329__i18__net5 n402__i18__net5 45
rk505 n336__i18__net5 n403__i18__net5 45
rk506 n478__r_out n479__r_out 8.6557
rk507 n479__r_out n480__r_out 1.541
rk508 n480__r_out n474__r_out 31.89e-3
rk510 n478__r_out n479__r_out 3.75
rk511 n478__r_out n480__r_out 3.75
rk512 n482__r_out n483__r_out 8.8496
rk513 n483__r_out n477__r_out 105.1e-3
rk514 n477__r_out n484__r_out 1.4342
rk515 n484__r_out n482__r_out 4.641
rk516 n482__r_out n483__r_out 3.1
rk517 n482__r_out n484__r_out 3.1
rk518 n339__i18__net5 n411__i18__net5 45.5
rk519 n346__i18__net5 n416__i18__net5 45
rk520 n493__r_out n494__r_out 8.6557
rk521 n494__r_out n495__r_out 1.541
rk522 n495__r_out n487__r_out 40.59e-3
rk524 n493__r_out n494__r_out 3.75
rk525 n493__r_out n495__r_out 3.75
rk526 n497__r_out n498__r_out 8.8496
rk527 n498__r_out n490__r_out 114.7e-3
rk528 n490__r_out n499__r_out 1.4246
rk529 n499__r_out n497__r_out 4.641
rk530 n497__r_out n498__r_out 3.1
rk531 n497__r_out n499__r_out 3.1
rk532 n349__i18__net5 n418__i18__net5 45.5
rk533 n1__x3 n2__x3 75.3305
rk534 n2__x3 n3__x3 62.2257
rk535 n1__x2 n2__x2 62.2257
rk536 n2__x2 n3__x2 75.3305
rk537 n1__x1 n2__x1 75.3305
rk538 n2__x1 n3__x1 62.2257
rk539 n1__x0 n2__x0 62.2257
rk540 n2__x0 n3__x0 75.3305
rk541 n8__ck n9__ck 4.733e-3
rk542 n10__ck n11__ck 4.733e-3
rk543 n9__ck n10__ck 12.55e-3
rk544 n2__ck n11__ck 45
rk545 n8__reset n9__reset 4.733e-3
rk546 n10__reset n11__reset 4.733e-3
rk547 n9__reset n10__reset 12.55e-3
rk548 n2__reset n11__reset 45
rk549 i14__net9 n17__i14__net9 509.5e-3
rk550 n18__i14__net9 n3__i14__net9 509.5e-3
rk551 n5__i14__net9 n19__i14__net9 509.5e-3
rk552 n20__i14__net9 n7__i14__net9 509.5e-3
rk553 n17__i14__net10 n18__i14__net10 3.427e-3
rk554 i14__net10 n19__i14__net10 3.427e-3
rk555 n17__i14__net10 n19__i14__net10 9.465e-3
rk556 n3__i14__net10 n20__i14__net10 3.427e-3
rk557 n21__i14__net10 n22__i14__net10 3.427e-3
rk558 n20__i14__net10 n21__i14__net10 9.465e-3
rk559 n23__i14__net10 n24__i14__net10 3.427e-3
rk560 n5__i14__net10 n25__i14__net10 3.427e-3
rk561 n23__i14__net10 n25__i14__net10 9.465e-3
rk562 n7__i14__net10 n26__i14__net10 3.427e-3
rk563 n27__i14__net10 n28__i14__net10 3.427e-3
rk564 n26__i14__net10 n27__i14__net10 9.465e-3
rk565 n5__i14__i17__net3 n6__i14__i17__net3 75.28
rk566 n6__i14__i17__net3 n7__i14__i17__net3 31.2971
rk567 n5__i14__i17__net6 n6__i14__i17__net6 31.4874
rk568 n6__i14__i17__net6 n7__i14__i17__net6 75.0874
rk569 n356__i18__net5 n426__i18__net5 45.5
rk570 n8__i14__i13__net1 n10__i14__i13__net1 75.3825
rk571 n10__i14__i13__net1 n11__i14__i13__net1 51.22e-3
rk572 n11__i14__i13__net1 n12__i14__i13__net1 62.2727
rk573 n11__i14__i13__net1 n13__i14__i13__net1 75.4286
rk574 n9__i14__i13__net1 n10__i14__i13__net1 62
rk575 n8__i14__i16__net1 n10__i14__i16__net1 75.3852
rk576 n10__i14__i16__net1 n11__i14__i16__net1 51.22e-3
rk577 n11__i14__i16__net1 n12__i14__i16__net1 75.4403
rk578 n11__i14__i16__net1 n13__i14__i16__net1 62.2858
rk579 n9__i14__i16__net1 n10__i14__i16__net1 62
rk580 n8__i14__i10__net1 n10__i14__i10__net1 75.3825
rk581 n10__i14__i10__net1 n11__i14__i10__net1 51.22e-3
rk582 n11__i14__i10__net1 n12__i14__i10__net1 62.2727
rk583 n11__i14__i10__net1 n13__i14__i10__net1 75.4286
rk584 n9__i14__i10__net1 n10__i14__i10__net1 62
rk585 n8__i14__i9__net1 n10__i14__i9__net1 75.3852
rk586 n10__i14__i9__net1 n11__i14__i9__net1 51.22e-3
rk587 n11__i14__i9__net1 n12__i14__i9__net1 75.4403
rk588 n11__i14__i9__net1 n13__i14__i9__net1 62.2858
rk589 n9__i14__i9__net1 n10__i14__i9__net1 62
rk590 n5__i14__i17__net1 n6__i14__i17__net1 75.3397
rk591 n6__i14__i17__net1 n7__i14__i17__net1 62.2257
rk592 i14__i17__net8 n2__i14__i17__net8 62.2257
rk593 n2__i14__i17__net8 n3__i14__i17__net8 75.3359
rk594 n506__r_out n507__r_out 8.6557
rk595 n507__r_out n508__r_out 1.541
rk596 n508__r_out n501__r_out 43.48e-3
rk598 n506__r_out n507__r_out 3.75
rk599 n506__r_out n508__r_out 3.75
rk600 n510__r_out n511__r_out 8.8496
rk601 n511__r_out n502__r_out 119.8e-3
rk602 n502__r_out n512__r_out 1.4232
rk603 n512__r_out n510__r_out 4.641
rk604 n510__r_out n511__r_out 3.1
rk605 n510__r_out n512__r_out 3.1
rk606 i14__i17__net3 n8__i14__i17__net3 509.5e-3
rk607 n10__i14__i17__net1 i14__i17__net1 509.5e-3
rk608 i14__i13__net2 n4__i14__i13__net2 45.8942
rk609 i14__i16__net2 n4__i14__i16__net2 45.8942
rk610 i14__i10__net2 n4__i14__i10__net2 45.8942
rk611 i14__i9__net2 n4__i14__i9__net2 45.8942
rk612 n12__ck n13__ck 3.427e-3
rk613 n4__ck n14__ck 3.427e-3
rk614 n12__ck n14__ck 9.465e-3
rk615 i14__i17__net7 n5__i14__i17__net7 3.427e-3
rk616 n6__i14__i17__net7 n7__i14__i17__net7 3.427e-3
rk617 n5__i14__i17__net7 n6__i14__i17__net7 9.465e-3
rk618 n361__i18__net5 n431__i18__net5 45.5
rk619 n8__i14__i17__i2__net1 n10__i14__i17__i2__net1 75.3825
rk620 n10__i14__i17__i2__net1 n11__i14__i17__i2__net1 51.22e-3
rk621 n11__i14__i17__i2__net1 n12__i14__i17__i2__net1 62.2727
rk622 n11__i14__i17__i2__net1 n13__i14__i17__i2__net1 75.4286
rk623 n9__i14__i17__i2__net1 n10__i14__i17__i2__net1 62
rk624 n8__i14__i17__i3__net1 n10__i14__i17__i3__net1 75.3852
rk625 n10__i14__i17__i3__net1 n11__i14__i17__i3__net1 51.22e-3
rk626 n11__i14__i17__i3__net1 n12__i14__i17__i3__net1 75.4403
rk627 n11__i14__i17__i3__net1 n13__i14__i17__i3__net1 62.2858
rk628 n9__i14__i17__i3__net1 n10__i14__i17__i3__net1 62
rk629 n366__i18__net5 n434__i18__net5 45
rk630 i14__i17__i2__net2 n4__i14__i17__i2__net2 45.8942
rk631 i14__i17__i3__net2 n4__i14__i17__i3__net2 45.8942
rk632 n49__i14__net10 n37__i14__net10 1.2059
rk633 n39__i14__net10 n50__i14__net10 1.2059
rk634 n51__i14__net10 n41__i14__net10 1.2059
rk635 n43__i14__net10 n52__i14__net10 1.2059
rk636 n517__r_out n518__r_out 8.6557
rk637 n518__r_out n519__r_out 1.541
rk638 n519__r_out n514__r_out 31.89e-3
rk640 n517__r_out n518__r_out 3.75
rk641 n517__r_out n519__r_out 3.75
rk642 n521__r_out n522__r_out 8.8496
rk643 n522__r_out n515__r_out 105.1e-3
rk644 n515__r_out n523__r_out 1.4342
rk645 n523__r_out n521__r_out 4.641
rk646 n521__r_out n522__r_out 3.1
rk647 n521__r_out n523__r_out 3.1
rk648 n41__i14__net9 n21__i14__net9 1.7109
rk649 n42__i14__net9 n23__i14__net9 1.7109
rk650 n43__i14__net9 n25__i14__net9 1.7109
rk651 n44__i14__net9 n27__i14__net9 1.7109
rk652 n369__i18__net5 n438__i18__net5 45.5
rk653 n14__i14__i13__net1 n15__i14__i13__net1 75.812
rk654 n14__i14__i16__net1 n15__i14__i16__net1 75.812
rk655 n14__i14__i10__net1 n15__i14__i10__net1 75.812
rk656 n14__i14__i9__net1 n15__i14__i9__net1 75.812
rk657 n21__i14__net3 i14__net3 4.237e-3
rk658 n10__i14__net3 n22__i14__net3 4.237e-3
rk659 n21__i14__net3 n22__i14__net3 23.66e-3
rk660 n11__i14__net3 n23__i14__net3 4.237e-3
rk661 n24__i14__net3 n3__i14__net3 4.237e-3
rk662 n23__i14__net3 n24__i14__net3 23.66e-3
rk663 n25__i14__net3 n5__i14__net3 4.237e-3
rk664 n14__i14__net3 n26__i14__net3 4.237e-3
rk665 n25__i14__net3 n26__i14__net3 23.66e-3
rk666 n15__i14__net3 n27__i14__net3 4.237e-3
rk667 n28__i14__net3 n7__i14__net3 4.237e-3
rk668 n27__i14__net3 n28__i14__net3 23.66e-3
rk669 n15__ck n16__ck 1.2059
rk670 n10__i14__i17__net7 n11__i14__i17__net7 1.2059
rk671 n376__i18__net5 n446__i18__net5 45
rk672 n10__i14__i17__net3 n9__i14__i17__net3 1.2109
rk673 n19__i14__i17__net1 n18__i14__i17__net1 1.2109
rk674 n526__r_out n527__r_out 8.6557
rk675 n527__r_out n528__r_out 1.541
rk676 n528__r_out n529__r_out 43.48e-3
rk678 n526__r_out n527__r_out 3.75
rk679 n526__r_out n528__r_out 3.75
rk680 n531__r_out n532__r_out 8.8496
rk681 n532__r_out n533__r_out 117.9e-3
rk682 n533__r_out n534__r_out 1.4214
rk683 n534__r_out n531__r_out 4.641
rk684 n531__r_out n532__r_out 3.1
rk685 n531__r_out n534__r_out 3.1
rk686 n4__i14__i13__net1 n16__i14__i13__net1 228.1e-3
rk687 n4__i14__i16__net1 n16__i14__i16__net1 228.1e-3
rk688 n4__i14__i10__net1 n16__i14__i10__net1 228.1e-3
rk689 n4__i14__i9__net1 n16__i14__i9__net1 228.1e-3
rk690 n14__i14__i17__i2__net1 n15__i14__i17__i2__net1 75.812
rk691 n14__i14__i17__i3__net1 n15__i14__i17__i3__net1 75.812
rk692 n16__reset n4__reset 4.237e-3
rk693 n17__reset n18__reset 4.237e-3
rk694 n16__reset n18__reset 23.66e-3
rk695 n19__reset n20__reset 4.237e-3
rk696 n21__reset n6__reset 4.237e-3
rk697 n20__reset n21__reset 23.66e-3
rk698 n379__i18__net5 n449__i18__net5 45
rk699 n4__i14__i17__i2__net1 n16__i14__i17__i2__net1 228.1e-3
rk700 n4__i14__i17__i3__net1 n16__i14__i17__i3__net1 228.1e-3
rk701 n386__i18__net5 n456__i18__net5 45
rk702 n6__i14__i13__net2 n7__i14__i13__net2 75.1559
rk703 n7__i14__i13__net2 n8__i14__i13__net2 277e-3
rk704 n8__i14__i13__net2 n10__i14__i13__net2 307.9e-3
rk705 n7__i14__i13__net2 n11__i14__i13__net2 62.4304
rk706 n8__i14__i13__net2 n12__i14__i13__net2 37.7116
rk707 n10__i14__i13__net2 n5__i14__i13__net2 108e-3
rk708 n9__i14__i13__net2 n10__i14__i13__net2 15.5
rk709 n6__i14__i16__net2 n7__i14__i16__net2 62.4304
rk710 n7__i14__i16__net2 n8__i14__i16__net2 277e-3
rk711 n8__i14__i16__net2 n9__i14__i16__net2 37.7116
rk712 n7__i14__i16__net2 n10__i14__i16__net2 75.1559
rk713 n8__i14__i16__net2 n12__i14__i16__net2 307.9e-3
rk714 n12__i14__i16__net2 n5__i14__i16__net2 112.8e-3
rk715 n11__i14__i16__net2 n12__i14__i16__net2 15.5
rk716 n6__i14__i10__net2 n7__i14__i10__net2 75.1559
rk717 n7__i14__i10__net2 n8__i14__i10__net2 277e-3
rk718 n8__i14__i10__net2 n10__i14__i10__net2 307.9e-3
rk719 n7__i14__i10__net2 n11__i14__i10__net2 62.4304
rk720 n8__i14__i10__net2 n12__i14__i10__net2 37.7116
rk721 n10__i14__i10__net2 n5__i14__i10__net2 108e-3
rk722 n9__i14__i10__net2 n10__i14__i10__net2 15.5
rk723 n6__i14__i9__net2 n7__i14__i9__net2 62.4304
rk724 n7__i14__i9__net2 n8__i14__i9__net2 277e-3
rk725 n8__i14__i9__net2 n9__i14__i9__net2 37.7116
rk726 n7__i14__i9__net2 n10__i14__i9__net2 75.1559
rk727 n8__i14__i9__net2 n12__i14__i9__net2 307.9e-3
rk728 n12__i14__i9__net2 n5__i14__i9__net2 112.8e-3
rk729 n11__i14__i9__net2 n12__i14__i9__net2 15.5
rk730 n539__r_out n540__r_out 8.6557
rk731 n540__r_out n541__r_out 1.541
rk732 n541__r_out n542__r_out 31.89e-3
rk734 n539__r_out n540__r_out 3.75
rk735 n539__r_out n541__r_out 3.75
rk736 n544__r_out n545__r_out 8.8496
rk737 n545__r_out n546__r_out 108.9e-3
rk738 n546__r_out n547__r_out 1.438
rk739 n547__r_out n544__r_out 4.641
rk740 n544__r_out n545__r_out 3.1
rk741 n544__r_out n547__r_out 3.1
rk742 n9__i14__net10 n53__i14__net10 509.5e-3
rk743 n9__i14__net9 n45__i14__net9 509.5e-3
rk744 n46__i14__net9 n11__i14__net9 509.5e-3
rk745 n54__i14__net10 n11__i14__net10 509.5e-3
rk746 n13__i14__net10 n55__i14__net10 509.5e-3
rk747 n13__i14__net9 n47__i14__net9 509.5e-3
rk748 n48__i14__net9 n15__i14__net9 509.5e-3
rk749 n56__i14__net10 n15__i14__net10 509.5e-3
rk750 n391__i18__net5 n461__i18__net5 45.5
rk751 n8__i14__i13__net5 n10__i14__i13__net5 75.3825
rk752 n10__i14__i13__net5 n11__i14__i13__net5 51.22e-3
rk753 n11__i14__i13__net5 n12__i14__i13__net5 62.2693
rk754 n11__i14__i13__net5 n13__i14__i13__net5 75.4286
rk755 n9__i14__i13__net5 n10__i14__i13__net5 62
rk756 n8__i14__i16__net5 n10__i14__i16__net5 75.3852
rk757 n10__i14__i16__net5 n11__i14__i16__net5 51.22e-3
rk758 n11__i14__i16__net5 n12__i14__i16__net5 75.4403
rk759 n11__i14__i16__net5 n13__i14__i16__net5 62.2822
rk760 n9__i14__i16__net5 n10__i14__i16__net5 62
rk761 n8__i14__i10__net5 n10__i14__i10__net5 75.3825
rk762 n10__i14__i10__net5 n11__i14__i10__net5 51.22e-3
rk763 n11__i14__i10__net5 n12__i14__i10__net5 62.2693
rk764 n11__i14__i10__net5 n13__i14__i10__net5 75.4286
rk765 n9__i14__i10__net5 n10__i14__i10__net5 62
rk766 n8__i14__i9__net5 n10__i14__i9__net5 75.3852
rk767 n10__i14__i9__net5 n11__i14__i9__net5 51.22e-3
rk768 n11__i14__i9__net5 n12__i14__i9__net5 75.4403
rk769 n11__i14__i9__net5 n13__i14__i9__net5 62.2822
rk770 n9__i14__i9__net5 n10__i14__i9__net5 62
rk771 n6__i14__i17__i2__net2 n7__i14__i17__i2__net2 75.1559
rk772 n7__i14__i17__i2__net2 n8__i14__i17__i2__net2 277e-3
rk773 n8__i14__i17__i2__net2 n10__i14__i17__i2__net2 307.9e-3
rk774 n7__i14__i17__i2__net2 n11__i14__i17__i2__net2 62.4304
rk775 n8__i14__i17__i2__net2 n12__i14__i17__i2__net2 37.7116
rk776 n10__i14__i17__i2__net2 n5__i14__i17__i2__net2 108e-3
rk777 n9__i14__i17__i2__net2 n10__i14__i17__i2__net2 15.5
rk778 n6__i14__i17__i3__net2 n7__i14__i17__i3__net2 62.4304
rk779 n7__i14__i17__i3__net2 n8__i14__i17__i3__net2 277e-3
rk780 n8__i14__i17__i3__net2 n9__i14__i17__i3__net2 37.7116
rk781 n7__i14__i17__i3__net2 n10__i14__i17__i3__net2 75.1559
rk782 n8__i14__i17__i3__net2 n12__i14__i17__i3__net2 307.9e-3
rk783 n12__i14__i17__i3__net2 n5__i14__i17__i3__net2 112.8e-3
rk784 n11__i14__i17__i3__net2 n12__i14__i17__i3__net2 15.5
rk785 n396__i18__net5 n467__i18__net5 45
rk786 n6__ck n21__ck 509.5e-3
rk787 n3__i14__i17__net3 n11__i14__i17__net3 509.5e-3
rk788 n20__i14__i17__net1 n3__i14__i17__net1 509.5e-3
rk789 n12__i14__i17__net7 n3__i14__i17__net7 509.5e-3
rk790 i14__i13__net4 n7__i14__i13__net4 45.8942
rk791 i14__i16__net4 n7__i14__i16__net4 45.8942
rk792 i14__i10__net4 n7__i14__i10__net4 45.8942
rk793 i14__i9__net4 n7__i14__i9__net4 45.8942
rk794 n552__r_out n553__r_out 8.6557
rk795 n553__r_out n554__r_out 1.541
rk796 n554__r_out n555__r_out 40.59e-3
rk798 n552__r_out n553__r_out 3.75
rk799 n552__r_out n554__r_out 3.75
rk800 n557__r_out n558__r_out 8.8496
rk801 n558__r_out n559__r_out 118.5e-3
rk802 n559__r_out n560__r_out 1.4283
rk803 n560__r_out n557__r_out 4.641
rk804 n557__r_out n558__r_out 3.1
rk805 n557__r_out n560__r_out 3.1
rk806 n399__i18__net5 n468__i18__net5 45.5
rk807 n8__i14__i17__i2__net5 n10__i14__i17__i2__net5 75.3825
rk808 n10__i14__i17__i2__net5 n11__i14__i17__i2__net5 51.22e-3
rk809 n11__i14__i17__i2__net5 n12__i14__i17__i2__net5 62.2693
rk810 n11__i14__i17__i2__net5 n13__i14__i17__i2__net5 75.4286
rk811 n9__i14__i17__i2__net5 n10__i14__i17__i2__net5 62
rk812 n8__i14__i17__i3__net5 n10__i14__i17__i3__net5 75.3852
rk813 n10__i14__i17__i3__net5 n11__i14__i17__i3__net5 51.22e-3
rk814 n11__i14__i17__i3__net5 n12__i14__i17__i3__net5 75.4403
rk815 n11__i14__i17__i3__net5 n13__i14__i17__i3__net5 62.2822
rk816 n9__i14__i17__i3__net5 n10__i14__i17__i3__net5 62
rk817 i14__i17__i2__net4 n7__i14__i17__i2__net4 45.8942
rk818 i14__i17__i3__net4 n7__i14__i17__i3__net4 45.8942
rk819 n2__i14__net4 n17__i14__net4 40.14e-3
rk820 n4__i14__net4 n18__i14__net4 40.14e-3
rk821 n6__i14__net4 n19__i14__net4 40.14e-3
rk822 n8__i14__net4 n20__i14__net4 40.14e-3
rk823 n406__i18__net5 n473__i18__net5 45.5
rk824 n565__r_out n566__r_out 8.6557
rk825 n566__r_out n567__r_out 1.541
rk826 n567__r_out n568__r_out 43.48e-3
rk828 n565__r_out n566__r_out 3.75
rk829 n565__r_out n567__r_out 3.75
rk830 n570__r_out n571__r_out 8.8496
rk831 n571__r_out n572__r_out 117.9e-3
rk832 n572__r_out n573__r_out 1.4214
rk833 n573__r_out n570__r_out 4.641
rk834 n570__r_out n571__r_out 3.1
rk835 n570__r_out n573__r_out 3.1
rk836 n4__i14__i13__net5 n14__i14__i13__net5 212e-3
rk837 n14__i14__i13__net5 n15__i14__i13__net5 62.0166
rk838 n4__i14__i16__net5 n14__i14__i16__net5 212e-3
rk839 n14__i14__i16__net5 n15__i14__i16__net5 62.0166
rk840 n4__i14__i10__net5 n14__i14__i10__net5 212e-3
rk841 n14__i14__i10__net5 n15__i14__i10__net5 62.0166
rk842 n4__i14__i9__net5 n14__i14__i9__net5 212e-3
rk843 n14__i14__i9__net5 n15__i14__i9__net5 62.0166
rk844 n409__i18__net5 n475__i18__net5 45.5
rk845 n2__i14__i17__net6 n10__i14__i17__net6 40.14e-3
rk846 n4__i14__i17__net6 n11__i14__i17__net6 40.14e-3
rk847 n8__i14__i13__net4 n9__i14__i13__net4 37.6937
rk848 n9__i14__i13__net4 n11__i14__i13__net4 290e-3
rk849 n11__i14__i13__net4 n12__i14__i13__net4 608e-3
rk850 n10__i14__i13__net4 n11__i14__i13__net4 15.5
rk851 n8__i14__i16__net4 n9__i14__i16__net4 37.6937
rk852 n9__i14__i16__net4 n11__i14__i16__net4 290e-3
rk853 n11__i14__i16__net4 n12__i14__i16__net4 612.8e-3
rk854 n10__i14__i16__net4 n11__i14__i16__net4 15.5
rk855 n8__i14__i10__net4 n9__i14__i10__net4 37.6937
rk856 n9__i14__i10__net4 n11__i14__i10__net4 290e-3
rk857 n11__i14__i10__net4 n12__i14__i10__net4 608e-3
rk858 n10__i14__i10__net4 n11__i14__i10__net4 15.5
rk859 n8__i14__i9__net4 n9__i14__i9__net4 37.6937
rk860 n9__i14__i9__net4 n11__i14__i9__net4 290e-3
rk861 n11__i14__i9__net4 n12__i14__i9__net4 612.8e-3
rk862 n10__i14__i9__net4 n11__i14__i9__net4 15.5
rk863 n414__i18__net5 n477__i18__net5 45.5
rk864 n4__i14__i17__i2__net5 n14__i14__i17__i2__net5 212e-3
rk865 n14__i14__i17__i2__net5 n15__i14__i17__i2__net5 62.0166
rk866 n4__i14__i17__i3__net5 n14__i14__i17__i3__net5 212e-3
rk867 n14__i14__i17__i3__net5 n15__i14__i17__i3__net5 62.0166
rk868 n578__r_out n579__r_out 8.6557
rk869 n579__r_out n580__r_out 1.541
rk870 n580__r_out n581__r_out 31.89e-3
rk872 n578__r_out n579__r_out 3.75
rk873 n578__r_out n580__r_out 3.75
rk874 n583__r_out n584__r_out 8.8496
rk875 n584__r_out n585__r_out 108.9e-3
rk876 n585__r_out n586__r_out 1.438
rk877 n586__r_out n583__r_out 4.641
rk878 n583__r_out n584__r_out 3.1
rk879 n583__r_out n586__r_out 3.1
rk880 n5__i14__i13__net4 n13__i14__i13__net4 45.5268
rk881 n5__i14__i16__net4 n13__i14__i16__net4 45.5268
rk882 n5__i14__i10__net4 n13__i14__i10__net4 45.5268
rk883 n5__i14__i9__net4 n13__i14__i9__net4 45.5268
rk884 n8__i14__i17__i2__net4 n9__i14__i17__i2__net4 37.6937
rk885 n9__i14__i17__i2__net4 n11__i14__i17__i2__net4 290e-3
rk886 n11__i14__i17__i2__net4 n12__i14__i17__i2__net4 608e-3
rk887 n10__i14__i17__i2__net4 n11__i14__i17__i2__net4 15.5
rk888 n8__i14__i17__i3__net4 n9__i14__i17__i3__net4 37.6937
rk889 n9__i14__i17__i3__net4 n11__i14__i17__i3__net4 290e-3
rk890 n11__i14__i17__i3__net4 n12__i14__i17__i3__net4 612.8e-3
rk891 n10__i14__i17__i3__net4 n11__i14__i17__i3__net4 15.5
rk892 n420__i18__net5 n479__i18__net5 45.5
rk893 n3__i14__y_out_b_3 n7__i14__y_out_b_3 119.8e-3
rk894 n7__i14__y_out_b_3 n8__i14__y_out_b_3 177e-3
rk895 n8__i14__y_out_b_3 n9__i14__y_out_b_3 15.5974
rk896 n7__i14__y_out_b_3 n10__i14__y_out_b_3 37.708
rk897 n3__i14__y_out_b_0 n7__i14__y_out_b_0 119.8e-3
rk898 n7__i14__y_out_b_0 n8__i14__y_out_b_0 37.708
rk899 n7__i14__y_out_b_0 n9__i14__y_out_b_0 177e-3
rk900 n9__i14__y_out_b_0 n10__i14__y_out_b_0 15.5974
rk901 n3__i14__x_out_b_2 n7__i14__x_out_b_2 119.8e-3
rk902 n7__i14__x_out_b_2 n8__i14__x_out_b_2 177e-3
rk903 n8__i14__x_out_b_2 n9__i14__x_out_b_2 15.5974
rk904 n7__i14__x_out_b_2 n10__i14__x_out_b_2 37.708
rk905 n3__i14__x_out_b_3 n7__i14__x_out_b_3 119.8e-3
rk906 n7__i14__x_out_b_3 n8__i14__x_out_b_3 37.708
rk907 n7__i14__x_out_b_3 n9__i14__x_out_b_3 177e-3
rk908 n9__i14__x_out_b_3 n10__i14__x_out_b_3 15.5974
rk909 n424__i18__net5 n481__i18__net5 45
rk910 n5__i14__i17__i2__net4 n13__i14__i17__i2__net4 45.0268
rk911 n5__i14__i17__i3__net4 n13__i14__i17__i3__net4 45.0268
rk912 n591__r_out n592__r_out 8.6557
rk913 n592__r_out n593__r_out 1.541
rk914 n593__r_out n594__r_out 40.59e-3
rk916 n591__r_out n592__r_out 3.75
rk917 n591__r_out n593__r_out 3.75
rk918 n596__r_out n597__r_out 8.8496
rk919 n597__r_out n598__r_out 119.8e-3
rk920 n598__r_out n599__r_out 1.4232
rk921 n599__r_out n596__r_out 4.641
rk922 n596__r_out n597__r_out 3.1
rk923 n596__r_out n599__r_out 3.1
rk924 x_out_3 n2__x_out_3 37.655
rk925 n2__x_out_3 n3__x_out_3 15.8098
rk926 x_out_2 n2__x_out_2 15.8098
rk927 n2__x_out_2 n3__x_out_2 37.655
rk928 x_out_1 n2__x_out_1 37.655
rk929 n2__x_out_1 n3__x_out_1 15.8098
rk930 x_out_0 n2__x_out_0 15.8098
rk931 n2__x_out_0 n3__x_out_0 37.655
rk932 n429__i18__net5 n483__i18__net5 45.5
rk933 n16__i14__i17__net1 n26__i14__i17__net1 119.8e-3
rk934 n26__i14__i17__net1 n27__i14__i17__net1 177e-3
rk935 n27__i14__i17__net1 n28__i14__i17__net1 15.5974
rk936 n26__i14__i17__net1 n29__i14__i17__net1 37.708
rk937 n8__i14__i17__net8 n19__i14__i17__net8 119.8e-3
rk938 n19__i14__i17__net8 n20__i14__i17__net8 37.708
rk939 n19__i14__i17__net8 n21__i14__i17__net8 177e-3
rk940 n21__i14__i17__net8 n22__i14__i17__net8 15.5974
rk941 n1__y3 n2__y3 75.3305
rk942 n2__y3 n3__y3 62.2257
rk943 n1__y2 n2__y2 62.2257
rk944 n2__y2 n3__y2 75.3305
rk945 n1__y1 n2__y1 75.3305
rk946 n2__y1 n3__y1 62.2257
rk947 n1__y0 n2__y0 62.2257
rk948 n2__y0 n3__y0 75.3305
rk949 n33__i14__net9 n57__i14__net9 509.5e-3
rk950 n58__i14__net9 n35__i14__net9 509.5e-3
rk951 n37__i14__net9 n59__i14__net9 509.5e-3
rk952 n60__i14__net9 n39__i14__net9 509.5e-3
rk953 n17__i14__i17__net7 n18__i14__i17__net7 37.655
rk954 n18__i14__i17__net7 n19__i14__i17__net7 15.8098
rk955 n10__i14__i17__net11 n11__i14__i17__net11 15.8098
rk956 n11__i14__i17__net11 n12__i14__i17__net11 37.655
rk957 n65__i14__net10 n66__i14__net10 3.427e-3
rk958 n29__i14__net10 n67__i14__net10 3.427e-3
rk959 n65__i14__net10 n67__i14__net10 9.465e-3
rk960 n31__i14__net10 n68__i14__net10 3.427e-3
rk961 n69__i14__net10 n70__i14__net10 3.427e-3
rk962 n68__i14__net10 n69__i14__net10 9.465e-3
rk963 n71__i14__net10 n72__i14__net10 3.427e-3
rk964 n33__i14__net10 n73__i14__net10 3.427e-3
rk965 n71__i14__net10 n73__i14__net10 9.465e-3
rk966 n35__i14__net10 n74__i14__net10 3.427e-3
rk967 n75__i14__net10 n76__i14__net10 3.427e-3
rk968 n74__i14__net10 n75__i14__net10 9.465e-3
rk969 n436__i18__net5 n485__i18__net5 45.5
rk970 n604__r_out n605__r_out 8.6557
rk971 n605__r_out n606__r_out 1.541
rk972 n606__r_out n607__r_out 28.99e-3
rk974 n604__r_out n605__r_out 3.75
rk975 n604__r_out n606__r_out 3.75
rk976 n609__r_out n610__r_out 8.8496
rk977 n610__r_out n611__r_out 105.1e-3
rk978 n611__r_out n612__r_out 1.4342
rk979 n612__r_out n609__r_out 4.641
rk980 n609__r_out n610__r_out 3.1
rk981 n609__r_out n612__r_out 3.1
rk982 n8__i14__i11__net1 n10__i14__i11__net1 75.3825
rk983 n10__i14__i11__net1 n11__i14__i11__net1 51.22e-3
rk984 n11__i14__i11__net1 n12__i14__i11__net1 62.2727
rk985 n11__i14__i11__net1 n13__i14__i11__net1 75.4286
rk986 n9__i14__i11__net1 n10__i14__i11__net1 62
rk987 n8__i14__i14__net1 n10__i14__i14__net1 75.3852
rk988 n10__i14__i14__net1 n11__i14__i14__net1 51.22e-3
rk989 n11__i14__i14__net1 n12__i14__i14__net1 75.4403
rk990 n11__i14__i14__net1 n13__i14__i14__net1 62.2858
rk991 n9__i14__i14__net1 n10__i14__i14__net1 62
rk992 n8__i14__i15__net1 n10__i14__i15__net1 75.3825
rk993 n10__i14__i15__net1 n11__i14__i15__net1 51.22e-3
rk994 n11__i14__i15__net1 n12__i14__i15__net1 62.2727
rk995 n11__i14__i15__net1 n13__i14__i15__net1 75.4286
rk996 n9__i14__i15__net1 n10__i14__i15__net1 62
rk997 n8__i14__i12__net1 n10__i14__i12__net1 75.3852
rk998 n10__i14__i12__net1 n11__i14__i12__net1 51.22e-3
rk999 n11__i14__i12__net1 n12__i14__i12__net1 75.4403
rk1000 n11__i14__i12__net1 n13__i14__i12__net1 62.2858
rk1001 n9__i14__i12__net1 n10__i14__i12__net1 62
rk1002 n441__i18__net5 n487__i18__net5 45
rk1003 n3__i14__i17__net10 n9__i14__i17__net10 1.714e-3
rk1004 n11__i14__i17__net8 n23__i14__i17__net8 505.7e-3
rk1005 i14__i11__net2 n4__i14__i11__net2 45.8942
rk1006 i14__i14__net2 n4__i14__i14__net2 45.8942
rk1007 i14__i15__net2 n4__i14__i15__net2 45.8942
rk1008 i14__i12__net2 n4__i14__i12__net2 45.8942
rk1009 n25__i14__net11 n27__i14__net11 37.988
rk1010 n27__i14__net11 n28__i14__net11 587.8e-3
rk1011 n26__i14__net11 n27__i14__net11 15.5
rk1012 n8__i14__i17__net9 n9__i14__i17__net9 31.3254
rk1013 n9__i14__i17__net9 n10__i14__i17__net9 75.0967
rk1014 n13__i14__i17__net11 i14__i17__net11 4.733e-3
rk1015 n444__i18__net5 n489__i18__net5 45.5
rk1016 n24__i14__i17__net8 n12__i14__i17__net8 1.3602
rk1017 n3__i14__i17__net9 n11__i14__i17__net9 1.714e-3
rk1018 n617__r_out n618__r_out 8.6557
rk1019 n618__r_out n619__r_out 1.541
rk1020 n619__r_out n620__r_out 37.69e-3
rk1022 n617__r_out n618__r_out 3.75
rk1023 n617__r_out n619__r_out 3.75
rk1024 n622__r_out n623__r_out 8.8496
rk1025 n623__r_out n624__r_out 114.7e-3
rk1026 n624__r_out n625__r_out 1.4246
rk1027 n625__r_out n622__r_out 4.641
rk1028 n622__r_out n623__r_out 3.1
rk1029 n622__r_out n625__r_out 3.1
rk1030 n25__i14__net7 n27__i14__net7 15.9844
rk1031 n27__i14__net7 n28__i14__net7 505.8e-3
rk1032 n26__i14__net7 n27__i14__net7 37.5
rk1033 n77__i14__net10 n78__i14__net10 1.2059
rk1034 n79__i14__net10 n80__i14__net10 1.2059
rk1035 n81__i14__net10 n82__i14__net10 1.2059
rk1036 n83__i14__net10 n84__i14__net10 1.2059
rk1037 n14__i14__i17__net9 n15__i14__i17__net9 3.878e-3
rk1038 n16__i14__i17__net9 n17__i14__i17__net9 3.878e-3
rk1039 n15__i14__i17__net9 n16__i14__i17__net9 16.56e-3
rk1040 n6__i14__i17__net9 n17__i14__i17__net9 45
rk1041 n451__i18__net5 n491__i18__net5 45.5
rk1042 n73__i14__net9 n61__i14__net9 1.7109
rk1043 n74__i14__net9 n63__i14__net9 1.7109
rk1044 n75__i14__net9 n65__i14__net9 1.7109
rk1045 n76__i14__net9 n67__i14__net9 1.7109
rk1046 n11__i14__i17__net10 n12__i14__i17__net10 15.7094
rk1047 n12__i14__i17__net10 n13__i14__i17__net10 37.7613
rk1048 n14__i14__i11__net1 n15__i14__i11__net1 75.812
rk1049 n14__i14__i14__net1 n15__i14__i14__net1 75.812
rk1050 n14__i14__i15__net1 n15__i14__i15__net1 75.812
rk1051 n14__i14__i12__net1 n15__i14__i12__net1 75.812
rk1052 n454__i18__net5 n493__i18__net5 45.5
rk1053 n18__i14__i17__net9 n19__i14__i17__net9 15.8469
rk1054 n19__i14__i17__net9 n20__i14__i17__net9 37.6238
rk1055 n49__i14__net4 n50__i14__net4 37.8495
rk1056 n50__i14__net4 n51__i14__net4 15.6319
rk1057 n37__i14__net3 n29__i14__net3 4.237e-3
rk1058 n38__i14__net3 n39__i14__net3 4.237e-3
rk1059 n37__i14__net3 n39__i14__net3 23.66e-3
rk1060 n40__i14__net3 n41__i14__net3 4.237e-3
rk1061 n42__i14__net3 n31__i14__net3 4.237e-3
rk1062 n41__i14__net3 n42__i14__net3 23.66e-3
rk1063 n43__i14__net3 n33__i14__net3 4.237e-3
rk1064 n44__i14__net3 n45__i14__net3 4.237e-3
rk1065 n43__i14__net3 n45__i14__net3 23.66e-3
rk1066 n46__i14__net3 n47__i14__net3 4.237e-3
rk1067 n48__i14__net3 n35__i14__net3 4.237e-3
rk1068 n47__i14__net3 n48__i14__net3 23.66e-3
rk1069 n630__r_out n631__r_out 8.6557
rk1070 n631__r_out n632__r_out 1.541
rk1071 n632__r_out n633__r_out 40.59e-3
rk1073 n630__r_out n631__r_out 3.75
rk1074 n630__r_out n632__r_out 3.75
rk1075 n635__r_out n636__r_out 8.8496
rk1076 n636__r_out n637__r_out 119.8e-3
rk1077 n637__r_out n638__r_out 1.4232
rk1078 n638__r_out n635__r_out 4.641
rk1079 n635__r_out n636__r_out 3.1
rk1080 n635__r_out n638__r_out 3.1
rk1081 n14__i14__i17__net10 n15__i14__i17__net10 3.878e-3
rk1082 n16__i14__i17__net10 n17__i14__i17__net10 3.878e-3
rk1083 n15__i14__i17__net10 n16__i14__i17__net10 16.56e-3
rk1084 n6__i14__i17__net10 n14__i14__i17__net10 45
rk1085 n32__reset n48__reset 45.5
rk1086 n4__i14__i11__net1 n16__i14__i11__net1 228.1e-3
rk1087 n4__i14__i14__net1 n16__i14__i14__net1 228.1e-3
rk1088 n4__i14__i15__net1 n16__i14__i15__net1 228.1e-3
rk1089 n4__i14__i12__net1 n16__i14__i12__net1 228.1e-3
rk1090 n459__i18__net5 n495__i18__net5 45
rk1091 n52__i14__net4 n53__i14__net4 37.8638
rk1092 n53__i14__net4 n54__i14__net4 15.6319
rk1093 n5__i14__i17__net11 n14__i14__i17__net11 1.4981
rk1094 n49__reset n29__reset 45.5017
rk1095 n25__i14__i17__net8 n16__i14__i17__net8 1.886e-3
rk1096 n464__i18__net5 n497__i18__net5 45
rk1097 n18__i14__i17__net10 n19__i14__i17__net10 31.181
rk1098 n19__i14__i17__net10 n20__i14__i17__net10 75.2412
rk1099 n55__i14__net4 n56__i14__net4 37.8495
rk1100 n56__i14__net4 n57__i14__net4 15.6319
rk1101 n7__i14__i17__net11 n15__i14__i17__net11 5.657e-3
rk1102 n643__r_out n644__r_out 8.6557
rk1103 n644__r_out n645__r_out 1.541
rk1104 n645__r_out n646__r_out 28.99e-3
rk1106 n643__r_out n644__r_out 3.75
rk1107 n643__r_out n645__r_out 3.75
rk1108 n648__r_out n649__r_out 8.8496
rk1109 n649__r_out n650__r_out 105.1e-3
rk1110 n650__r_out n651__r_out 1.4342
rk1111 n651__r_out n648__r_out 4.641
rk1112 n648__r_out n649__r_out 3.1
rk1113 n648__r_out n651__r_out 3.1
rk1114 n6__i14__i11__net2 n7__i14__i11__net2 75.1559
rk1115 n7__i14__i11__net2 n8__i14__i11__net2 271.7e-3
rk1116 n8__i14__i11__net2 n10__i14__i11__net2 307.9e-3
rk1117 n7__i14__i11__net2 n11__i14__i11__net2 62.4304
rk1118 n8__i14__i11__net2 n12__i14__i11__net2 37.7116
rk1119 n10__i14__i11__net2 n5__i14__i11__net2 108e-3
rk1120 n9__i14__i11__net2 n10__i14__i11__net2 15.5
rk1121 n6__i14__i14__net2 n7__i14__i14__net2 62.4304
rk1122 n7__i14__i14__net2 n8__i14__i14__net2 277e-3
rk1123 n8__i14__i14__net2 n9__i14__i14__net2 37.7116
rk1124 n7__i14__i14__net2 n10__i14__i14__net2 75.1559
rk1125 n8__i14__i14__net2 n12__i14__i14__net2 307.9e-3
rk1126 n12__i14__i14__net2 n5__i14__i14__net2 112.8e-3
rk1127 n11__i14__i14__net2 n12__i14__i14__net2 15.5
rk1128 n6__i14__i15__net2 n7__i14__i15__net2 75.1559
rk1129 n7__i14__i15__net2 n8__i14__i15__net2 277e-3
rk1130 n8__i14__i15__net2 n10__i14__i15__net2 307.9e-3
rk1131 n7__i14__i15__net2 n11__i14__i15__net2 62.4304
rk1132 n8__i14__i15__net2 n12__i14__i15__net2 37.7116
rk1133 n10__i14__i15__net2 n5__i14__i15__net2 108e-3
rk1134 n9__i14__i15__net2 n10__i14__i15__net2 15.5
rk1135 n6__i14__i12__net2 n7__i14__i12__net2 62.4304
rk1136 n7__i14__i12__net2 n8__i14__i12__net2 277e-3
rk1137 n8__i14__i12__net2 n9__i14__i12__net2 37.7116
rk1138 n7__i14__i12__net2 n10__i14__i12__net2 75.1559
rk1139 n8__i14__i12__net2 n12__i14__i12__net2 307.9e-3
rk1140 n12__i14__i12__net2 n5__i14__i12__net2 112.8e-3
rk1141 n11__i14__i12__net2 n12__i14__i12__net2 15.5
rk1142 n471__i18__net5 n499__i18__net5 22.625
rk1143 n57__i14__net10 n93__i14__net10 509.5e-3
rk1144 n49__i14__net9 n77__i14__net9 509.5e-3
rk1145 n78__i14__net9 n51__i14__net9 509.5e-3
rk1146 n94__i14__net10 n59__i14__net10 509.5e-3
rk1147 n61__i14__net10 n95__i14__net10 509.5e-3
rk1148 n53__i14__net9 n79__i14__net9 509.5e-3
rk1149 n80__i14__net9 n55__i14__net9 509.5e-3
rk1150 n96__i14__net10 n63__i14__net10 509.5e-3
rk1151 n57__i14__net3 n58__i14__net3 15.9159
rk1152 n58__i14__net3 n59__i14__net3 37.5
rk1153 n8__i14__i11__net5 n10__i14__i11__net5 75.3825
rk1154 n10__i14__i11__net5 n11__i14__i11__net5 51.22e-3
rk1155 n11__i14__i11__net5 n12__i14__i11__net5 62.2693
rk1156 n11__i14__i11__net5 n13__i14__i11__net5 75.4286
rk1157 n9__i14__i11__net5 n10__i14__i11__net5 62
rk1158 n8__i14__i14__net5 n10__i14__i14__net5 75.3852
rk1159 n10__i14__i14__net5 n11__i14__i14__net5 51.22e-3
rk1160 n11__i14__i14__net5 n12__i14__i14__net5 75.4403
rk1161 n11__i14__i14__net5 n13__i14__i14__net5 62.2822
rk1162 n9__i14__i14__net5 n10__i14__i14__net5 62
rk1163 n8__i14__i15__net5 n10__i14__i15__net5 75.3825
rk1164 n10__i14__i15__net5 n11__i14__i15__net5 51.22e-3
rk1165 n11__i14__i15__net5 n12__i14__i15__net5 62.2693
rk1166 n11__i14__i15__net5 n13__i14__i15__net5 75.4286
rk1167 n9__i14__i15__net5 n10__i14__i15__net5 62
rk1168 n8__i14__i12__net5 n10__i14__i12__net5 75.3852
rk1169 n10__i14__i12__net5 n11__i14__i12__net5 51.22e-3
rk1170 n11__i14__i12__net5 n12__i14__i12__net5 75.4403
rk1171 n11__i14__i12__net5 n13__i14__i12__net5 62.2822
rk1172 n9__i14__i12__net5 n10__i14__i12__net5 62
rk1173 n70__i14__net4 n35__i14__net4 45.5017
rk1174 n3__i14__net7 n33__i14__net7 26.85e-3
rk1175 n33__i14__net7 n29__i14__net7 174.7e-3
rk1176 i14__i11__net4 n7__i14__i11__net4 45.8942
rk1177 i14__i14__net4 n7__i14__i14__net4 45.8942
rk1178 i14__i15__net4 n7__i14__i15__net4 45.8942
rk1179 i14__i12__net4 n7__i14__i12__net4 45.8942
rk1180 n60__i14__net3 n61__i14__net3 15.9302
rk1181 n61__i14__net3 n62__i14__net3 37.5
rk1182 i14__clk_div4_out_b n3__i14__clk_div4_out_b 16.014
rk1184 n2__i14__clk_div4_out_b n3__i14__clk_div4_out_b 37.5
rk1185 n32__i14__net4 n71__i14__net4 45.5
rk1186 n70__i14__net3 n68__i14__net3 15.9159
rk1187 n68__i14__net3 n71__i14__net3 37.5
rk1188 n22__i14__net4 n72__i14__net4 40.14e-3
rk1189 n24__i14__net4 n73__i14__net4 40.14e-3
rk1190 n26__i14__net4 n74__i14__net4 40.14e-3
rk1191 n28__i14__net4 n75__i14__net4 40.14e-3
rk1192 n3__i14__net11 n31__i14__net11 374.8e-3
rk1193 ck4 n3__ck4 37.9709
rk1194 n3__ck4 n4__ck4 583.1e-3
rk1195 n2__ck4 n3__ck4 15.5
rk1196 n4__i14__i11__net5 n14__i14__i11__net5 212e-3
rk1197 n14__i14__i11__net5 n15__i14__i11__net5 62.0166
rk1198 n4__i14__i14__net5 n14__i14__i14__net5 212e-3
rk1199 n14__i14__i14__net5 n15__i14__i14__net5 62.0166
rk1200 n4__i14__i15__net5 n14__i14__i15__net5 212e-3
rk1201 n14__i14__i15__net5 n15__i14__i15__net5 62.0166
rk1202 n4__i14__i12__net5 n14__i14__i12__net5 212e-3
rk1203 n14__i14__i12__net5 n15__i14__i12__net5 62.0166
rk1204 n9__i14__i11__net4 n10__i14__i11__net4 37.6937
rk1205 n10__i14__i11__net4 n12__i14__i11__net4 290e-3
rk1206 n12__i14__i11__net4 n8__i14__i11__net4 108e-3
rk1207 n11__i14__i11__net4 n12__i14__i11__net4 15.5
rk1208 n9__i14__i14__net4 n10__i14__i14__net4 37.6937
rk1209 n10__i14__i14__net4 n12__i14__i14__net4 290e-3
rk1210 n12__i14__i14__net4 n8__i14__i14__net4 112.8e-3
rk1211 n11__i14__i14__net4 n12__i14__i14__net4 15.5
rk1212 n9__i14__i15__net4 n10__i14__i15__net4 37.6937
rk1213 n10__i14__i15__net4 n12__i14__i15__net4 290e-3
rk1214 n12__i14__i15__net4 n8__i14__i15__net4 108e-3
rk1215 n11__i14__i15__net4 n12__i14__i15__net4 15.5
rk1216 n9__i14__i12__net4 n10__i14__i12__net4 37.6937
rk1217 n10__i14__i12__net4 n12__i14__i12__net4 290e-3
rk1218 n12__i14__i12__net4 n8__i14__i12__net4 112.8e-3
rk1219 n11__i14__i12__net4 n12__i14__i12__net4 15.5
rk1220 n86__i14__net9 n87__i14__net9 37.8463
rk1221 n87__i14__net9 n88__i14__net9 15.6359
rk1222 n97__i14__net10 n98__i14__net10 15.9159
rk1223 n98__i14__net10 n99__i14__net10 37.5
rk1224 n2__i18__net4 n43__i18__net4 45
rk1225 n11__i14__net7 n34__i14__net7 45
rk1226 n11__i14__net11 n34__i14__net11 45
rk1227 n506__i18__net5 n507__i18__net5 13.5129
rk1228 n507__i18__net5 n508__i18__net5 1.541
rk1229 n508__i18__net5 n502__i18__net5 46.38e-3
rk1231 n506__i18__net5 n507__i18__net5 3.75
rk1232 n506__i18__net5 n508__i18__net5 3.75
rk1233 n510__i18__net5 n511__i18__net5 16.4166
rk1234 n511__i18__net5 n505__i18__net5 463.3e-3
rk1235 n505__i18__net5 n512__i18__net5 1.0573
rk1236 n512__i18__net5 n510__i18__net5 4.641
rk1237 n510__i18__net5 n511__i18__net5 3.2632
rk1238 n510__i18__net5 n512__i18__net5 3.1
rk1239 n89__i14__net9 n90__i14__net9 37.8606
rk1240 n90__i14__net9 n91__i14__net9 15.6359
rk1241 n100__i14__net10 n101__i14__net10 15.9302
rk1242 n101__i14__net10 n102__i14__net10 37.5
rk1243 n5__i14__i11__net4 n13__i14__i11__net4 45.0268
rk1244 n5__i14__i14__net4 n13__i14__i14__net4 45.0268
rk1245 n5__i14__i15__net4 n13__i14__i15__net4 45.0268
rk1246 n5__i14__i12__net4 n13__i14__i12__net4 45.0268
rk1247 n5__i18__net4 n51__i18__net4 45.5
rk1248 n8__i14__net7 n37__i14__net7 45.5
rk1249 n8__i14__net11 n36__i14__net11 45.5
rk1250 n8__i18__net4 n56__i18__net4 45.5
rk1251 n92__i14__net9 n93__i14__net9 37.8463
rk1252 n93__i14__net9 n94__i14__net9 15.6359
rk1253 n103__i14__net10 n104__i14__net10 15.9159
rk1254 n104__i14__net10 n105__i14__net10 37.5
rk1255 n3__i14__x_out_b_1 n7__i14__x_out_b_1 119.8e-3
rk1256 n7__i14__x_out_b_1 n8__i14__x_out_b_1 177e-3
rk1257 n8__i14__x_out_b_1 n9__i14__x_out_b_1 15.5974
rk1258 n7__i14__x_out_b_1 n10__i14__x_out_b_1 37.708
rk1259 n3__i14__y_out_b_2 n7__i14__y_out_b_2 119.8e-3
rk1260 n7__i14__y_out_b_2 n8__i14__y_out_b_2 37.708
rk1261 n7__i14__y_out_b_2 n9__i14__y_out_b_2 177e-3
rk1262 n9__i14__y_out_b_2 n10__i14__y_out_b_2 15.5974
rk1263 n3__i14__y_out_b_1 n7__i14__y_out_b_1 119.8e-3
rk1264 n7__i14__y_out_b_1 n8__i14__y_out_b_1 177e-3
rk1265 n8__i14__y_out_b_1 n9__i14__y_out_b_1 15.5974
rk1266 n7__i14__y_out_b_1 n10__i14__y_out_b_1 37.708
rk1267 n3__i14__x_out_b_0 n7__i14__x_out_b_0 119.8e-3
rk1268 n7__i14__x_out_b_0 n8__i14__x_out_b_0 37.708
rk1269 n7__i14__x_out_b_0 n9__i14__x_out_b_0 177e-3
rk1270 n9__i14__x_out_b_0 n10__i14__x_out_b_0 15.5974
rk1271 n515__i18__net5 n516__i18__net5 13.5129
rk1272 n516__i18__net5 n517__i18__net5 1.541
rk1273 n517__i18__net5 n518__i18__net5 34.79e-3
rk1275 n515__i18__net5 n516__i18__net5 3.75
rk1276 n515__i18__net5 n517__i18__net5 3.75
rk1277 n520__i18__net5 n521__i18__net5 16.4166
rk1278 n521__i18__net5 n522__i18__net5 450.5e-3
rk1279 n522__i18__net5 n523__i18__net5 1.0701
rk1280 n523__i18__net5 n520__i18__net5 4.641
rk1281 n520__i18__net5 n521__i18__net5 3.2632
rk1282 n520__i18__net5 n523__i18__net5 3.1
rk1283 n7__y_out_3 n8__y_out_3 37.655
rk1284 n8__y_out_3 n9__y_out_3 15.8098
rk1285 n7__y_out_2 n8__y_out_2 15.8098
rk1286 n8__y_out_2 n9__y_out_2 37.655
rk1287 n7__y_out_1 n8__y_out_1 37.655
rk1288 n8__y_out_1 n9__y_out_1 15.8098
rk1289 n9__y_out_0 n10__y_out_0 15.8098
rk1290 n10__y_out_0 n11__y_out_0 37.655
rk1291 n11__i18__net4 n58__i18__net4 45.5
rk1292 n5__ck_b n6__ck_b 37.8274
rk1293 n6__ck_b n7__ck_b 15.643
rk1294 n14__i18__net4 n66__i18__net4 45
rk1295 n8__x_out_2 n16__x_out_2 6.854e-3
rk1296 n3__y_out_0 n14__y_out_0 6.854e-3
rk1297 n528__i18__net5 n529__i18__net5 13.5129
rk1298 n529__i18__net5 n530__i18__net5 1.541
rk1299 n530__i18__net5 n531__i18__net5 43.48e-3
rk1301 n528__i18__net5 n529__i18__net5 3.75
rk1302 n528__i18__net5 n530__i18__net5 3.75
rk1303 n533__i18__net5 n534__i18__net5 16.4166
rk1304 n534__i18__net5 n535__i18__net5 460.1e-3
rk1305 n535__i18__net5 n536__i18__net5 1.0605
rk1306 n536__i18__net5 n533__i18__net5 4.641
rk1307 n533__i18__net5 n534__i18__net5 3.2632
rk1308 n533__i18__net5 n536__i18__net5 3.1
rk1309 n3__i13__i14__net2 n4__i13__i14__net2 75.0403
rk1310 n4__i13__i14__net2 n5__i13__i14__net2 31.3601
rk1311 n3__i13__i12__net2 n4__i13__i12__net2 31.3601
rk1312 n4__i13__i12__net2 n5__i13__i12__net2 75.0403
rk1313 n11__net11 n4__net11 45.5171
rk1314 n6__ck4 n7__ck4 62.2257
rk1315 n7__ck4 n8__ck4 75.3305
rk1316 n17__i18__net4 n71__i18__net4 45.5
rk1317 n8__ck_b ck_b 509.5e-3
rk1318 n9__ck_b n10__ck_b 37.8349
rk1319 n10__ck_b n11__ck_b 15.66
rk1320 ck_buff n5__ck_buff 3.427e-3
rk1321 n6__ck_buff n7__ck_buff 3.427e-3
rk1322 n5__ck_buff n6__ck_buff 9.465e-3
rk1323 n12__y_out_2 n13__y_out_2 75.4527
rk1324 n13__y_out_2 n14__y_out_2 62.0153
rk1325 n14__x_out_0 n15__x_out_0 75.4527
rk1326 n15__x_out_0 n16__x_out_0 62.0153
rk1327 n11__x_out_2 n21__x_out_2 55.48e-3
rk1328 n21__x_out_2 n17__x_out_2 490.2e-3
rk1329 n6__y_out_0 n17__y_out_0 55.48e-3
rk1330 n17__y_out_0 n15__y_out_0 490.2e-3
rk1331 n6__i13__i14__net2 n2__i13__i14__net2 3.514e-3
rk1332 n2__i13__i12__net2 n6__i13__i12__net2 3.514e-3
rk1333 n8__i9__i4__net1 n10__i9__i4__net1 75.3852
rk1334 n10__i9__i4__net1 n11__i9__i4__net1 51.22e-3
rk1335 n11__i9__i4__net1 n12__i9__i4__net1 75.4403
rk1336 n11__i9__i4__net1 n13__i9__i4__net1 62.2858
rk1337 n9__i9__i4__net1 n10__i9__i4__net1 62
rk1338 n9__i13__a2 n11__i13__a2 75.4649
rk1339 n11__i13__a2 n12__i13__a2 519.5e-3
rk1340 n10__i13__a2 n11__i13__a2 62
rk1341 n9__i13__a0 n11__i13__a0 75.4649
rk1342 n11__i13__a0 n12__i13__a0 519.9e-3
rk1343 n10__i13__a0 n11__i13__a0 62
rk1344 n20__i18__net4 n76__i18__net4 45
rk1345 n541__i18__net5 n542__i18__net5 13.5129
rk1346 n542__i18__net5 n543__i18__net5 1.541
rk1347 n543__i18__net5 n544__i18__net5 46.38e-3
rk1349 n541__i18__net5 n542__i18__net5 3.75
rk1350 n541__i18__net5 n543__i18__net5 3.75
rk1351 n546__i18__net5 n547__i18__net5 16.4166
rk1352 n547__i18__net5 n548__i18__net5 463.3e-3
rk1353 n548__i18__net5 n549__i18__net5 1.0573
rk1354 n549__i18__net5 n546__i18__net5 4.641
rk1355 n546__i18__net5 n547__i18__net5 3.2632
rk1356 n546__i18__net5 n549__i18__net5 3.1
rk1357 i9__i4__net2 n4__i9__i4__net2 45.8942
rk1358 n22__x_out_2 n23__x_out_2 31.6782
rk1359 n18__y_out_0 n19__y_out_0 31.6782
rk1360 n7__i13__i14__net2 n8__i13__i14__net2 6.35e-3
rk1361 n9__i13__i14__net2 n11__i13__i14__net2 6.35e-3
rk1362 n8__i13__i14__net2 n9__i13__i14__net2 28.4e-3
rk1363 n10__i13__i14__net2 n11__i13__i14__net2 75
rk1364 n7__i13__i12__net2 n9__i13__i12__net2 6.35e-3
rk1365 n10__i13__i12__net2 n11__i13__i12__net2 6.35e-3
rk1366 n7__i13__i12__net2 n11__i13__i12__net2 28.4e-3
rk1367 n8__i13__i12__net2 n9__i13__i12__net2 75
rk1368 n3__y_out_2 n19__y_out_2 212.1e-3
rk1369 n8__x_out_0 n19__x_out_0 212.1e-3
rk1370 n23__i18__net4 n78__i18__net4 45.5
rk1371 n15__i13__a2 n17__i13__a2 75.3453
rk1372 n17__i13__a2 n18__i13__a2 561.7e-3
rk1373 n16__i13__a2 n17__i13__a2 31
rk1374 n16__i13__a0 n17__i13__a0 561.7e-3
rk1375 n16__i13__a0 n18__i13__a0 75.3453
rk1376 n15__i13__a0 n16__i13__a0 31
rk1377 n13__net11 n14__net11 75.1706
rk1378 n14__net11 n15__net11 184.8e-3
rk1379 n15__net11 n12__net11 189.4e-3
rk1380 n12__net11 net11 17.08e-3
rk1381 n14__net11 n16__net11 31.2187
rk1382 n15__net11 n17__net11 31.2044
rk1383 n15__net11 n18__net11 75.1616
rk1384 n10__ck_buff n11__ck_buff 1.2059
rk1385 n26__i18__net4 n86__i18__net4 45.5
rk1386 n560__i18__net5 n561__i18__net5 13.5129
rk1387 n561__i18__net5 n562__i18__net5 1.541
rk1388 n562__i18__net5 n554__i18__net5 34.79e-3
rk1390 n560__i18__net5 n561__i18__net5 3.75
rk1391 n560__i18__net5 n562__i18__net5 3.75
rk1392 n564__i18__net5 n565__i18__net5 16.4166
rk1393 n565__i18__net5 n557__i18__net5 450.5e-3
rk1394 n557__i18__net5 n566__i18__net5 1.0701
rk1395 n566__i18__net5 n564__i18__net5 4.641
rk1396 n564__i18__net5 n565__i18__net5 3.2632
rk1397 n564__i18__net5 n566__i18__net5 3.1
rk1398 n17__ck_b n16__ck_b 1.2109
rk1399 n14__i9__i4__net1 n15__i9__i4__net1 75.812
rk1400 n29__i18__net4 n91__i18__net4 45
rk1401 n3__reset_buff n4__reset_buff 4.237e-3
rk1402 n5__reset_buff reset_buff 4.237e-3
rk1403 n4__reset_buff n5__reset_buff 23.66e-3
rk1404 n32__i18__net4 n94__i18__net4 45
rk1405 n4__i9__i4__net1 n16__i9__i4__net1 228.1e-3
rk1406 n8__x_out_3 n17__x_out_3 6.854e-3
rk1407 n8__x_out_1 n16__x_out_1 6.854e-3
rk1408 n11__net9 n12__net9 75.1652
rk1409 n12__net9 net9 305.3e-3
rk1410 n12__net9 n13__net9 31.208
rk1411 n567__i18__net5 n568__i18__net5 13.5129
rk1412 n568__i18__net5 n569__i18__net5 1.541
rk1413 n569__i18__net5 n570__i18__net5 46.38e-3
rk1415 n567__i18__net5 n568__i18__net5 3.75
rk1416 n567__i18__net5 n569__i18__net5 3.75
rk1417 n572__i18__net5 n573__i18__net5 16.4166
rk1418 n573__i18__net5 n574__i18__net5 463.3e-3
rk1419 n574__i18__net5 n575__i18__net5 1.0573
rk1420 n575__i18__net5 n572__i18__net5 4.641
rk1421 n572__i18__net5 n573__i18__net5 3.2632
rk1422 n572__i18__net5 n575__i18__net5 3.1
rk1423 n3__i13__i15__net2 n4__i13__i15__net2 75.0403
rk1424 n4__i13__i15__net2 n5__i13__i15__net2 31.3601
rk1425 n3__i13__i13__net2 n4__i13__i13__net2 31.3601
rk1426 n4__i13__i13__net2 n5__i13__i13__net2 75.0403
rk1427 n35__i18__net4 n98__i18__net4 45.5
rk1428 n7__reset_b n8__reset_b 37.8274
rk1429 n8__reset_b n9__reset_b 15.643
rk1430 n30__ck n22__ck 524.4e-3
rk1431 n13__y_out_3 n14__y_out_3 75.4527
rk1432 n14__y_out_3 n15__y_out_3 62.0153
rk1433 n12__y_out_1 n13__y_out_1 75.4527
rk1434 n13__y_out_1 n14__y_out_1 62.0153
rk1435 n11__x_out_3 n20__x_out_3 55.48e-3
rk1436 n20__x_out_3 n18__x_out_3 490.2e-3
rk1437 n11__x_out_1 n19__x_out_1 55.48e-3
rk1438 n19__x_out_1 n17__x_out_1 490.2e-3
rk1439 n6__i13__i15__net2 n2__i13__i15__net2 3.514e-3
rk1440 n2__i13__i13__net2 n6__i13__i13__net2 3.514e-3
rk1441 n11__net12 n4__net12 45.5171
rk1442 n6__i9__i4__net2 n7__i9__i4__net2 62.4304
rk1443 n7__i9__i4__net2 n8__i9__i4__net2 277e-3
rk1444 n8__i9__i4__net2 n9__i9__i4__net2 37.7116
rk1445 n7__i9__i4__net2 n10__i9__i4__net2 75.1559
rk1446 n8__i9__i4__net2 n12__i9__i4__net2 307.9e-3
rk1447 n12__i9__i4__net2 n5__i9__i4__net2 112.8e-3
rk1448 n11__i9__i4__net2 n12__i9__i4__net2 15.5
rk1449 n38__i18__net4 n106__i18__net4 45.5
rk1450 n9__i13__a3 n11__i13__a3 75.4649
rk1451 n11__i13__a3 n12__i13__a3 519.5e-3
rk1452 n10__i13__a3 n11__i13__a3 62
rk1453 n9__i13__a1 n11__i13__a1 75.4649
rk1454 n11__i13__a1 n12__i13__a1 519.9e-3
rk1455 n10__i13__a1 n11__i13__a1 62
rk1456 n10__reset_b n11__reset_b 37.8349
rk1457 n11__reset_b n12__reset_b 15.66
rk1458 n580__i18__net5 n581__i18__net5 13.5129
rk1459 n581__i18__net5 n582__i18__net5 1.541
rk1460 n582__i18__net5 n583__i18__net5 34.79e-3
rk1462 n580__i18__net5 n581__i18__net5 3.75
rk1463 n580__i18__net5 n582__i18__net5 3.75
rk1464 n585__i18__net5 n586__i18__net5 16.4166
rk1465 n586__i18__net5 n587__i18__net5 448.6e-3
rk1466 n587__i18__net5 n588__i18__net5 1.0682
rk1467 n588__i18__net5 n585__i18__net5 4.641
rk1468 n585__i18__net5 n586__i18__net5 3.2632
rk1469 n585__i18__net5 n588__i18__net5 3.1
rk1470 n18__ck_b n3__ck_b 509.5e-3
rk1471 n12__ck_buff n3__ck_buff 509.5e-3
rk1472 n21__x_out_3 n22__x_out_3 31.6782
rk1473 n22__x_out_1 n23__x_out_1 31.6782
rk1474 n7__i13__i15__net2 n8__i13__i15__net2 6.35e-3
rk1475 n9__i13__i15__net2 n11__i13__i15__net2 6.35e-3
rk1476 n8__i13__i15__net2 n9__i13__i15__net2 28.4e-3
rk1477 n10__i13__i15__net2 n11__i13__i15__net2 75
rk1478 n7__i13__i13__net2 n9__i13__i13__net2 6.35e-3
rk1479 n10__i13__i13__net2 n11__i13__i13__net2 6.35e-3
rk1480 n7__i13__i13__net2 n11__i13__i13__net2 28.4e-3
rk1481 n8__i13__i13__net2 n9__i13__i13__net2 75
rk1482 n3__y_out_3 n18__y_out_3 212.1e-3
rk1483 n3__y_out_1 n19__y_out_1 212.1e-3
rk1484 n41__i18__net4 n108__i18__net4 45.5
rk1485 n8__i9__i4__net5 n10__i9__i4__net5 75.3852
rk1486 n10__i9__i4__net5 n11__i9__i4__net5 51.22e-3
rk1487 n11__i9__i4__net5 n12__i9__i4__net5 75.4403
rk1488 n11__i9__i4__net5 n13__i9__i4__net5 62.2822
rk1489 n9__i9__i4__net5 n10__i9__i4__net5 62
rk1490 n13__i13__a3 n15__i13__a3 75.3453
rk1491 n15__i13__a3 n16__i13__a3 561.7e-3
rk1492 n14__i13__a3 n15__i13__a3 31
rk1493 n14__i13__a1 n15__i13__a1 561.7e-3
rk1494 n14__i13__a1 n16__i13__a1 75.3453
rk1495 n13__i13__a1 n14__i13__a1 31
rk1496 i9__i4__net4 n7__i9__i4__net4 45.8942
rk1497 n46__i18__net4 n116__i18__net4 45.5
rk1498 n599__i18__net5 n600__i18__net5 13.5129
rk1499 n600__i18__net5 n601__i18__net5 1.541
rk1500 n601__i18__net5 n593__i18__net5 43.48e-3
rk1502 n599__i18__net5 n600__i18__net5 3.75
rk1503 n599__i18__net5 n601__i18__net5 3.75
rk1504 n603__i18__net5 n604__i18__net5 16.4166
rk1505 n604__i18__net5 n596__i18__net5 458.2e-3
rk1506 n596__i18__net5 n605__i18__net5 1.0586
rk1507 n605__i18__net5 n603__i18__net5 4.641
rk1508 n603__i18__net5 n604__i18__net5 3.2632
rk1509 n603__i18__net5 n605__i18__net5 3.1
rk1510 n13__net12 n14__net12 75.1706
rk1511 n14__net12 n15__net12 184.8e-3
rk1512 n15__net12 n12__net12 172.3e-3
rk1513 n12__net12 net12 17.08e-3
rk1514 n14__net12 n16__net12 31.2187
rk1515 n15__net12 n17__net12 31.2044
rk1516 n15__net12 n18__net12 75.1616
rk1517 n49__i18__net4 n119__i18__net4 45
rk1518 n2__reset_b n14__reset_b 40.14e-3
rk1519 n54__i18__net4 n123__i18__net4 45.5
rk1520 n5__i13__i17__net1 n6__i13__i17__net1 31.5319
rk1521 n5__i13__i16__net1 n6__i13__i16__net1 31.5319
rk1522 n3__i13__a3 n19__i13__a3 513.2e-3
rk1523 n3__i13__a1 n19__i13__a1 513.2e-3
rk1524 n4__i9__i4__net5 n14__i9__i4__net5 212e-3
rk1525 n14__i9__i4__net5 n15__i9__i4__net5 62.0166
rk1526 n606__i18__net5 n607__i18__net5 13.5129
rk1527 n607__i18__net5 n608__i18__net5 1.541
rk1528 n608__i18__net5 n609__i18__net5 46.38e-3
rk1530 n606__i18__net5 n607__i18__net5 3.75
rk1531 n606__i18__net5 n608__i18__net5 3.75
rk1532 n611__i18__net5 n612__i18__net5 16.4166
rk1533 n612__i18__net5 n613__i18__net5 463.3e-3
rk1534 n613__i18__net5 n614__i18__net5 1.0573
rk1535 n614__i18__net5 n611__i18__net5 4.641
rk1536 n611__i18__net5 n612__i18__net5 3.2632
rk1537 n611__i18__net5 n614__i18__net5 3.1
rk1538 n11__net10 n12__net10 75.1652
rk1539 n12__net10 net10 180.9e-3
rk1540 n12__net10 n13__net10 31.208
rk1541 n28__ck n34__ck 195.6e-3
rk1542 n3__i13__a2 n23__i13__a2 511.3e-3
rk1543 n3__i13__a0 n23__i13__a0 511.3e-3
rk1544 n60__i18__net4 n125__i18__net4 45.5
rk1545 n8__i9__i4__net4 n9__i9__i4__net4 37.6937
rk1546 n9__i9__i4__net4 n11__i9__i4__net4 290e-3
rk1547 n11__i9__i4__net4 n12__i9__i4__net4 612.8e-3
rk1548 n10__i9__i4__net4 n11__i9__i4__net4 15.5
rk1549 n51__reset n60__reset 338.7e-3
rk1550 n64__i18__net4 n127__i18__net4 45.5
rk1551 n8__i13__i17__net1 n9__i13__i17__net1 37.7009
rk1552 n9__i13__i17__net1 n7__i13__i17__net1 283.1e-3
rk1553 n7__i13__i17__net1 n10__i13__i17__net1 31
rk1554 n9__i13__i17__net1 n3__i13__i17__net1 170.8e-3
rk1555 n8__i13__i16__net1 n9__i13__i16__net1 37.7009
rk1556 n9__i13__i16__net1 n7__i13__i16__net1 282.9e-3
rk1557 n7__i13__i16__net1 n10__i13__i16__net1 31
rk1558 n9__i13__i16__net1 n3__i13__i16__net1 170.8e-3
rk1559 n9__net13 n11__net13 17.08e-3
rk1560 n11__net13 n12__net13 163.8e-3
rk1561 n12__net13 n13__net13 31.208
rk1562 n12__net13 n14__net13 75.1652
rk1563 n5__i9__i4__net4 n13__i9__i4__net4 45.5268
rk1564 n619__i18__net5 n620__i18__net5 13.5129
rk1565 n620__i18__net5 n621__i18__net5 1.541
rk1566 n621__i18__net5 n622__i18__net5 34.79e-3
rk1568 n619__i18__net5 n620__i18__net5 3.75
rk1569 n619__i18__net5 n621__i18__net5 3.75
rk1570 n624__i18__net5 n625__i18__net5 16.4166
rk1571 n625__i18__net5 n626__i18__net5 448.6e-3
rk1572 n626__i18__net5 n627__i18__net5 1.0682
rk1573 n627__i18__net5 n624__i18__net5 4.641
rk1574 n624__i18__net5 n625__i18__net5 3.2632
rk1575 n624__i18__net5 n627__i18__net5 3.1
rk1576 n13__ck_buff n14__ck_buff 37.8349
rk1577 n14__ck_buff n15__ck_buff 15.66
rk1578 n57__reset n63__reset 285.5e-3
rk1579 n9__i13__net11 n11__i13__net11 554.6e-3
rk1580 n11__i13__net11 n12__i13__net11 31.3424
rk1581 n10__i13__net11 n11__i13__net11 75
rk1582 n11__i13__net1 n13__i13__net1 554.6e-3
rk1583 n13__i13__net1 n14__i13__net1 31.3424
rk1584 n12__i13__net1 n13__i13__net1 75
rk1585 n69__i18__net4 n129__i18__net4 45
rk1586 n2__net13 n15__net13 45.0171
rk1587 n3__i9__net2 n5__i9__net2 119.8e-3
rk1588 n5__i9__net2 n6__i9__net2 37.708
rk1589 n5__i9__net2 n7__i9__net2 177e-3
rk1590 n7__i9__net2 n8__i9__net2 15.5974
rk1591 n7__i13__a2 n24__i13__a2 6.854e-3
rk1592 n7__i13__a0 n24__i13__a0 6.854e-3
rk1593 n24__ck_buff n25__ck_buff 37.8274
rk1594 n25__ck_buff n26__ck_buff 15.643
rk1595 n74__i18__net4 n131__i18__net4 45.5
rk1596 n7__i9__net1 n8__i9__net1 15.8098
rk1597 n8__i9__net1 n9__i9__net1 37.655
rk1598 n3__i13__i17__i4__net2 n4__i13__i17__i4__net2 75.0403
rk1599 n4__i13__i17__i4__net2 n5__i13__i17__i4__net2 31.3601
rk1600 n3__i13__i16__i4__net2 n4__i13__i16__i4__net2 31.3601
rk1601 n4__i13__i16__i4__net2 n5__i13__i16__i4__net2 75.0403
rk1602 n11__net14 n12__net14 75.1632
rk1603 n12__net14 n13__net14 31.2096
rk1604 n12__net14 n14__net14 165.9e-3
rk1605 n14__net14 n9__net14 17.08e-3
rk1606 n638__i18__net5 n639__i18__net5 13.5129
rk1607 n639__i18__net5 n640__i18__net5 1.541
rk1608 n640__i18__net5 n636__i18__net5 43.48e-3
rk1610 n638__i18__net5 n639__i18__net5 3.75
rk1611 n638__i18__net5 n640__i18__net5 3.75
rk1612 n642__i18__net5 n643__i18__net5 16.4166
rk1613 n643__i18__net5 n637__i18__net5 463.3e-3
rk1614 n637__i18__net5 n644__i18__net5 1.0573
rk1615 n644__i18__net5 n642__i18__net5 4.641
rk1616 n642__i18__net5 n643__i18__net5 3.2632
rk1617 n642__i18__net5 n644__i18__net5 3.1
rk1618 n10__reset_buff n11__reset_buff 37.8349
rk1619 n11__reset_buff n12__reset_buff 15.66
rk1620 n20__i13__a3 n21__i13__a3 75.4527
rk1621 n21__i13__a3 n22__i13__a3 62.0153
rk1622 n20__i13__a1 n21__i13__a1 75.4527
rk1623 n21__i13__a1 n22__i13__a1 62.0153
rk1624 n81__i18__net4 n133__i18__net4 45.5
rk1625 n14__i13__a2 n27__i13__a2 55.48e-3
rk1626 n27__i13__a2 n25__i13__a2 490.2e-3
rk1627 n14__i13__a0 n27__i13__a0 55.48e-3
rk1628 n27__i13__a0 n25__i13__a0 490.2e-3
rk1629 n6__i13__i17__i4__net2 n2__i13__i17__i4__net2 3.514e-3
rk1630 n2__i13__i16__i4__net2 n6__i13__i16__i4__net2 3.514e-3
rk1631 i9__i1__net1 n2__i9__i1__net1 25.5752
rk1632 n2__net14 n15__net14 45.5171
rk1633 n9__i13__net12 n11__i13__net12 75.4649
rk1634 n11__i13__net12 n12__i13__net12 519.5e-3
rk1635 n10__i13__net12 n11__i13__net12 62
rk1636 n11__i13__net2 n13__i13__net2 75.4649
rk1637 n13__i13__net2 n14__i13__net2 519.9e-3
rk1638 n12__i13__net2 n13__i13__net2 62
rk1639 n3__i9__net1 n10__i9__net1 45.0568
rk1640 n25__shift n26__shift 21.2464
rk1641 n27__shift n28__shift 25.5797
rk1642 n84__i18__net4 n135__i18__net4 45.5
rk1643 n13__reset_buff n14__reset_buff 37.8274
rk1644 n14__reset_buff n15__reset_buff 15.643
rk1645 n28__i13__a2 n29__i13__a2 31.6782
rk1646 n28__i13__a0 n29__i13__a0 31.6782
rk1647 n7__i13__i17__i4__net2 n8__i13__i17__i4__net2 6.35e-3
rk1648 n9__i13__i17__i4__net2 n11__i13__i17__i4__net2 6.35e-3
rk1649 n8__i13__i17__i4__net2 n9__i13__i17__i4__net2 28.4e-3
rk1650 n10__i13__i17__i4__net2 n11__i13__i17__i4__net2 75
rk1651 n7__i13__i16__i4__net2 n9__i13__i16__i4__net2 6.35e-3
rk1652 n10__i13__i16__i4__net2 n11__i13__i16__i4__net2 6.35e-3
rk1653 n7__i13__i16__i4__net2 n11__i13__i16__i4__net2 28.4e-3
rk1654 n8__i13__i16__i4__net2 n9__i13__i16__i4__net2 75
rk1655 n645__i18__net5 n646__i18__net5 13.5129
rk1656 n646__i18__net5 n647__i18__net5 1.541
rk1657 n647__i18__net5 n648__i18__net5 31.89e-3
rk1659 n645__i18__net5 n646__i18__net5 3.75
rk1660 n645__i18__net5 n647__i18__net5 3.75
rk1661 n650__i18__net5 n651__i18__net5 16.4166
rk1662 n651__i18__net5 n652__i18__net5 450.5e-3
rk1663 n652__i18__net5 n653__i18__net5 1.0701
rk1664 n653__i18__net5 n650__i18__net5 4.641
rk1665 n650__i18__net5 n651__i18__net5 3.2632
rk1666 n650__i18__net5 n653__i18__net5 3.1
rk1667 n7__i13__a3 n24__i13__a3 212.1e-3
rk1668 n7__i13__a1 n24__i13__a1 212.1e-3
rk1669 n3__i9__i1__net1 n4__i9__i1__net1 25.5797
rk1670 n13__i13__net12 n15__i13__net12 75.3453
rk1671 n15__i13__net12 n16__i13__net12 561.7e-3
rk1672 n14__i13__net12 n15__i13__net12 31
rk1673 n16__i13__net2 n17__i13__net2 561.7e-3
rk1674 n16__i13__net2 n18__i13__net2 75.3453
rk1675 n15__i13__net2 n16__i13__net2 31
rk1676 n89__i18__net4 n137__i18__net4 45.5
rk1677 n12__ck4 n16__ck4 45.0502
rk1678 n29__shift n30__shift 21.2464
rk1679 n6__i9__i1__net1 n5__i9__i1__net1 25.0752
rk1680 n96__i18__net4 n139__i18__net4 45.5
rk1681 n658__i18__net5 n659__i18__net5 13.5129
rk1682 n659__i18__net5 n660__i18__net5 1.541
rk1683 n660__i18__net5 n661__i18__net5 40.59e-3
rk1685 n658__i18__net5 n659__i18__net5 3.75
rk1686 n658__i18__net5 n660__i18__net5 3.75
rk1687 n663__i18__net5 n664__i18__net5 16.4166
rk1688 n664__i18__net5 n665__i18__net5 460.1e-3
rk1689 n665__i18__net5 n666__i18__net5 1.0605
rk1690 n666__i18__net5 n663__i18__net5 4.641
rk1691 n663__i18__net5 n664__i18__net5 3.2632
rk1692 n663__i18__net5 n666__i18__net5 3.1
rk1693 n101__i18__net4 n141__i18__net4 45.5
rk1694 n31__shift n3__shift 2.521e-3
rk1695 n32__shift n7__shift 2.521e-3
rk1696 n33__shift n11__shift 2.521e-3
rk1697 n5__i2__net79 n7__i2__net79 550.1e-3
rk1698 n7__i2__net79 n8__i2__net79 342.8e-3
rk1699 n8__i2__net79 n9__i2__net79 31.1609
rk1700 n6__i2__net79 n7__i2__net79 75
rk1701 n5__i1__net79 n7__i1__net79 550.1e-3
rk1702 n7__i1__net79 n8__i1__net79 342.8e-3
rk1703 n8__i1__net79 n9__i1__net79 31.1609
rk1704 n6__i1__net79 n7__i1__net79 75
rk1705 n5__i0__net79 n7__i0__net79 550.1e-3
rk1706 n7__i0__net79 n8__i0__net79 342.8e-3
rk1707 n8__i0__net79 n9__i0__net79 31.1609
rk1708 n6__i0__net79 n7__i0__net79 75
rk1709 n5__i13__i19__net1 n6__i13__i19__net1 31.5319
rk1710 n5__i13__i18__net1 n6__i13__i18__net1 31.5319
rk1711 n3__i13__net11 n15__i13__net11 513.2e-3
rk1712 n3__i13__net12 n19__i13__net12 513.2e-3
rk1713 n104__i18__net4 n143__i18__net4 45.5
rk1714 n4__net4 n2__net4 31.1339
rk1715 n2__net4 n5__net4 75.4173
rk1716 n4__net3 net3 31.1339
rk1717 net3 n5__net3 75.4173
rk1718 n528__vss n527__vss 31.1339
rk1719 n527__vss n529__vss 75.4173
rk1720 n10__i2__net79 n2__i2__net79 3.134e-3
rk1721 n10__i1__net79 n2__i1__net79 3.134e-3
rk1722 n10__i0__net79 n2__i0__net79 3.134e-3
rk1723 n677__i18__net5 n678__i18__net5 13.5129
rk1724 n678__i18__net5 n679__i18__net5 1.541
rk1725 n679__i18__net5 n672__i18__net5 43.48e-3
rk1727 n677__i18__net5 n678__i18__net5 3.75
rk1728 n677__i18__net5 n679__i18__net5 3.75
rk1729 n681__i18__net5 n682__i18__net5 16.4166
rk1730 n682__i18__net5 n673__i18__net5 463.3e-3
rk1731 n673__i18__net5 n683__i18__net5 1.0573
rk1732 n683__i18__net5 n681__i18__net5 4.641
rk1733 n681__i18__net5 n682__i18__net5 3.2632
rk1734 n681__i18__net5 n683__i18__net5 3.1
rk1735 n3__i13__net1 n17__i13__net1 511.3e-3
rk1736 n3__i13__net2 n21__i13__net2 511.3e-3
rk1737 n14__shift n34__shift 3.001e-3
rk1738 n35__shift n16__shift 3.001e-3
rk1739 n18__shift n36__shift 3.001e-3
rk1740 n111__i18__net4 n145__i18__net4 45.5
rk1741 n11__i2__net79 n4__i2__net79 503.2e-3
rk1742 n11__i1__net79 n4__i1__net79 503.2e-3
rk1743 n11__i0__net79 n4__i0__net79 503.2e-3
rk1744 n37__shift n19__shift 2.751e-3
rk1745 n21__shift n38__shift 2.751e-3
rk1746 n39__shift n23__shift 2.751e-3
rk1747 n3__r0_buff n4__r0_buff 31.0977
rk1748 n4__r0_buff n5__r0_buff 75.3952
rk1749 n3__r1_buff n4__r1_buff 31.0977
rk1750 n4__r1_buff n5__r1_buff 75.3952
rk1751 n3__r2_buff n4__r2_buff 31.0977
rk1752 n4__r2_buff n5__r2_buff 75.3952
rk1753 n8__i13__i19__net1 n9__i13__i19__net1 37.7009
rk1754 n9__i13__i19__net1 n7__i13__i19__net1 283.1e-3
rk1755 n7__i13__i19__net1 n10__i13__i19__net1 31
rk1756 n9__i13__i19__net1 n3__i13__i19__net1 170.8e-3
rk1757 n8__i13__i18__net1 n9__i13__i18__net1 37.7009
rk1758 n9__i13__i18__net1 n7__i13__i18__net1 282.9e-3
rk1759 n7__i13__i18__net1 n10__i13__i18__net1 31
rk1760 n9__i13__i18__net1 n3__i13__i18__net1 170.8e-3
rk1761 n114__i18__net4 n147__i18__net4 45.5
rk1762 n5__i13__net17 n7__i13__net17 554.6e-3
rk1763 n7__i13__net17 n8__i13__net17 31.3424
rk1764 n6__i13__net17 n7__i13__net17 75
rk1765 n9__i13__net7 n11__i13__net7 554.6e-3
rk1766 n11__i13__net7 n12__i13__net7 31.3424
rk1767 n10__i13__net7 n11__i13__net7 75
rk1768 n684__i18__net5 n685__i18__net5 13.5129
rk1769 n685__i18__net5 n686__i18__net5 1.541
rk1770 n686__i18__net5 n687__i18__net5 31.89e-3
rk1772 n684__i18__net5 n685__i18__net5 3.75
rk1773 n684__i18__net5 n686__i18__net5 3.75
rk1774 n689__i18__net5 n690__i18__net5 16.4166
rk1775 n690__i18__net5 n691__i18__net5 450.5e-3
rk1776 n691__i18__net5 n692__i18__net5 1.0701
rk1777 n692__i18__net5 n689__i18__net5 4.641
rk1778 n689__i18__net5 n690__i18__net5 3.2632
rk1779 n689__i18__net5 n692__i18__net5 3.1
rk1780 n121__i18__net4 n149__i18__net4 22.625
rk1781 n7__i13__net1 n18__i13__net1 6.854e-3
rk1782 n7__i13__net2 n22__i13__net2 6.854e-3
rk1783 n535__vss n536__vss 4.2431
rk1784 n536__vss n537__vss 934.9e-3
rk1785 n537__vss n538__vss 72.47e-3
rk1786 n538__vss n539__vss 856e-3
rk1787 n539__vss n540__vss 129e-3
rk1788 n540__vss n541__vss 661.3e-3
rk1789 n541__vss n543__vss 334.1e-3
rk1790 n543__vss n532__vss 129e-3
rk1791 n532__vss n544__vss 856e-3
rk1792 n544__vss n533__vss 72.47e-3
rk1793 n533__vss n534__vss 934.9e-3
rk1794 n534__vss n542__vss 4.2431
rk1795 n541__vss n545__vss 174.4e-3
rk1796 n545__vss n546__vss 155.5e-3
rk1797 n546__vss n548__vss 334.1e-3
rk1798 n548__vss n523__vss 108.6e-3
rk1799 n523__vss n549__vss 856.6e-3
rk1800 n549__vss n524__vss 61.01e-3
rk1801 n524__vss n525__vss 924.1e-3
rk1802 n525__vss n547__vss 4.2377
rk1803 n546__vss n550__vss 329.9e-3
rk1804 n550__vss n552__vss 334.1e-3
rk1805 n552__vss n520__vss 108.6e-3
rk1806 n520__vss n553__vss 856.6e-3
rk1807 n553__vss n521__vss 61.01e-3
rk1808 n521__vss n522__vss 924.1e-3
rk1809 n522__vss n551__vss 4.2377
rk1810 n550__vss n554__vss 329.9e-3
rk1811 n554__vss n556__vss 334.1e-3
rk1812 n556__vss n517__vss 108.6e-3
rk1813 n517__vss n557__vss 856.6e-3
rk1814 n557__vss n518__vss 61.01e-3
rk1815 n518__vss n519__vss 924.1e-3
rk1816 n519__vss n555__vss 4.2377
rk1817 n554__vss n558__vss 329.9e-3
rk1818 n558__vss n560__vss 334.1e-3
rk1819 n560__vss n514__vss 108.6e-3
rk1820 n514__vss n561__vss 856.6e-3
rk1821 n561__vss n515__vss 61.01e-3
rk1822 n515__vss n516__vss 924.1e-3
rk1823 n516__vss n559__vss 4.2377
rk1824 n558__vss n562__vss 41.89e-3
rk1825 n562__vss n563__vss 288e-3
rk1826 n563__vss n565__vss 334.1e-3
rk1827 n565__vss n511__vss 118.8e-3
rk1828 n511__vss n566__vss 855.3e-3
rk1829 n566__vss n512__vss 66.71e-3
rk1830 n512__vss n513__vss 928.4e-3
rk1831 n513__vss n564__vss 4.2399
rk1832 n563__vss n567__vss 329.9e-3
rk1833 n567__vss n569__vss 334.1e-3
rk1834 n569__vss n500__vss 118.8e-3
rk1835 n500__vss n570__vss 855.3e-3
rk1836 n570__vss n501__vss 66.71e-3
rk1837 n501__vss n502__vss 928.4e-3
rk1838 n502__vss n568__vss 4.2399
rk1839 n567__vss n571__vss 329.9e-3
rk1840 n571__vss n573__vss 334.1e-3
rk1841 n573__vss n497__vss 93.21e-3
rk1842 n497__vss n574__vss 847.4e-3
rk1843 n574__vss n498__vss 52.36e-3
rk1844 n498__vss n575__vss 1.0029
rk1845 n575__vss n572__vss 4.3255
rk1846 n571__vss n576__vss 329.9e-3
rk1847 n576__vss n578__vss 334.1e-3
rk1848 n578__vss n494__vss 93.21e-3
rk1849 n494__vss n579__vss 847.4e-3
rk1850 n579__vss n495__vss 52.36e-3
rk1851 n495__vss n580__vss 1.0029
rk1852 n580__vss n577__vss 4.3255
rk1854 n576__vss n581__vss 41.89e-3
rk1855 n581__vss n582__vss 288e-3
rk1856 n582__vss n584__vss 334.1e-3
rk1857 n584__vss n491__vss 110.8e-3
rk1858 n491__vss n585__vss 856.6e-3
rk1859 n585__vss n492__vss 62.26e-3
rk1860 n492__vss n493__vss 925.3e-3
rk1861 n493__vss n583__vss 4.2383
rk1863 n582__vss n586__vss 329.9e-3
rk1864 n586__vss n588__vss 334.1e-3
rk1865 n588__vss n488__vss 118.8e-3
rk1866 n488__vss n589__vss 855.3e-3
rk1867 n589__vss n489__vss 66.71e-3
rk1868 n489__vss n490__vss 928.4e-3
rk1869 n490__vss n587__vss 4.2399
rk1870 n586__vss n590__vss 329.9e-3
rk1871 n590__vss n592__vss 334.1e-3
rk1872 n592__vss n485__vss 118.8e-3
rk1873 n485__vss n593__vss 855.3e-3
rk1874 n593__vss n486__vss 66.71e-3
rk1875 n486__vss n487__vss 928.4e-3
rk1876 n487__vss n591__vss 4.2399
rk1877 n590__vss n594__vss 329.9e-3
rk1878 n594__vss n596__vss 334.1e-3
rk1879 n596__vss n482__vss 120.4e-3
rk1880 n482__vss n597__vss 854.5e-3
rk1881 n597__vss n483__vss 67.65e-3
rk1882 n483__vss n484__vss 928.6e-3
rk1883 n484__vss n595__vss 4.24
rk1884 n594__vss n598__vss 41.89e-3
rk1885 n598__vss n599__vss 288e-3
rk1886 n599__vss n601__vss 334.1e-3
rk1887 n601__vss n479__vss 120.4e-3
rk1888 n479__vss n602__vss 854.5e-3
rk1889 n602__vss n480__vss 67.65e-3
rk1890 n480__vss n481__vss 928.6e-3
rk1891 n481__vss n600__vss 4.24
rk1892 n599__vss n604__vss 659.8e-3
rk1893 n604__vss n449__vss 129e-3
rk1894 n449__vss n605__vss 856e-3
rk1895 n605__vss n450__vss 72.47e-3
rk1896 n450__vss n451__vss 934.9e-3
rk1897 n451__vss n603__vss 4.2431
rk1898 n535__vss n538__vss 3.75
rk1899 n535__vss n540__vss 12.5
rk1900 n542__vss n543__vss 12.5
rk1901 n542__vss n544__vss 3.75
rk1902 n547__vss n548__vss 12.5
rk1903 n547__vss n549__vss 3.75
rk1904 n551__vss n552__vss 12.5
rk1905 n551__vss n553__vss 3.75
rk1906 n555__vss n556__vss 12.5
rk1907 n555__vss n557__vss 3.75
rk1908 n559__vss n560__vss 12.5
rk1909 n559__vss n561__vss 3.75
rk1910 n564__vss n565__vss 12.5
rk1911 n564__vss n566__vss 3.75
rk1912 n568__vss n569__vss 12.5
rk1913 n568__vss n570__vss 3.75
rk1914 n572__vss n573__vss 12.5
rk1915 n572__vss n574__vss 3.75
rk1916 n577__vss n578__vss 12.5
rk1917 n577__vss n579__vss 3.75
rk1918 n583__vss n584__vss 12.5
rk1919 n583__vss n585__vss 3.75
rk1920 n587__vss n588__vss 12.5
rk1921 n587__vss n589__vss 3.75
rk1922 n591__vss n592__vss 12.5
rk1923 n591__vss n593__vss 3.75
rk1924 n595__vss n596__vss 12.5
rk1925 n595__vss n597__vss 3.75
rk1926 n600__vss n601__vss 12.5
rk1927 n600__vss n602__vss 3.75
rk1928 n603__vss n604__vss 12.5
rk1929 n603__vss n605__vss 3.75
rk1930 n535__vddio n536__vddio 16.4166
rk1931 n536__vddio n537__vddio 769.2e-3
rk1932 n537__vddio n538__vddio 733.9e-3
rk1933 n538__vddio n539__vddio 560.6e-3
rk1934 n539__vddio n540__vddio 958.6e-3
rk1935 n540__vddio n541__vddio 213.8e-3
rk1936 n541__vddio n542__vddio 937.8e-3
rk1937 n542__vddio n543__vddio 174.4e-3
rk1938 n543__vddio n544__vddio 155.5e-3
rk1939 n544__vddio n545__vddio 329.9e-3
rk1940 n545__vddio n546__vddio 329.9e-3
rk1941 n546__vddio n547__vddio 329.9e-3
rk1942 n547__vddio n548__vddio 41.89e-3
rk1943 n548__vddio n549__vddio 288e-3
rk1944 n549__vddio n550__vddio 329.9e-3
rk1945 n550__vddio n551__vddio 329.9e-3
rk1946 n551__vddio n552__vddio 329.9e-3
rk1947 n552__vddio n553__vddio 41.89e-3
rk1948 n553__vddio n554__vddio 288e-3
rk1949 n554__vddio n555__vddio 329.9e-3
rk1950 n555__vddio n556__vddio 329.9e-3
rk1951 n556__vddio n557__vddio 329.9e-3
rk1952 n557__vddio n558__vddio 41.89e-3
rk1953 n558__vddio n559__vddio 288e-3
rk1954 n559__vddio n433__vddio 936.2e-3
rk1955 n542__vddio n533__vddio 610.5e-3
rk1956 n533__vddio n561__vddio 213.8e-3
rk1957 n561__vddio n532__vddio 958.6e-3
rk1958 n532__vddio n562__vddio 560.6e-3
rk1959 n562__vddio n529__vddio 733.9e-3
rk1960 n529__vddio n563__vddio 769.2e-3
rk1961 n563__vddio n560__vddio 16.4166
rk1962 n544__vddio n527__vddio 605.1e-3
rk1963 n527__vddio n565__vddio 208.4e-3
rk1964 n565__vddio n526__vddio 953.2e-3
rk1965 n526__vddio n566__vddio 555.1e-3
rk1966 n566__vddio n523__vddio 728.5e-3
rk1967 n523__vddio n567__vddio 763.8e-3
rk1968 n567__vddio n564__vddio 16.4166
rk1969 n545__vddio n521__vddio 605.1e-3
rk1970 n521__vddio n569__vddio 208.4e-3
rk1971 n569__vddio n520__vddio 953.2e-3
rk1972 n520__vddio n570__vddio 555.1e-3
rk1973 n570__vddio n517__vddio 728.5e-3
rk1974 n517__vddio n571__vddio 763.8e-3
rk1975 n571__vddio n568__vddio 16.4166
rk1976 n546__vddio n515__vddio 605.1e-3
rk1977 n515__vddio n573__vddio 208.4e-3
rk1978 n573__vddio n514__vddio 953.2e-3
rk1979 n514__vddio n574__vddio 555.1e-3
rk1980 n574__vddio n511__vddio 728.5e-3
rk1981 n511__vddio n575__vddio 763.8e-3
rk1982 n575__vddio n572__vddio 16.4166
rk1983 n547__vddio n510__vddio 605.1e-3
rk1984 n510__vddio n577__vddio 208.4e-3
rk1985 n577__vddio n507__vddio 953.2e-3
rk1986 n507__vddio n578__vddio 555.1e-3
rk1987 n578__vddio n506__vddio 728.5e-3
rk1988 n506__vddio n579__vddio 763.8e-3
rk1989 n579__vddio n576__vddio 16.4166
rk1990 n549__vddio n504__vddio 607.3e-3
rk1991 n504__vddio n581__vddio 210.6e-3
rk1992 n581__vddio n501__vddio 955.4e-3
rk1993 n501__vddio n582__vddio 557.3e-3
rk1994 n582__vddio n500__vddio 730.7e-3
rk1995 n500__vddio n583__vddio 766e-3
rk1996 n583__vddio n580__vddio 16.4166
rk1997 n550__vddio n497__vddio 607.3e-3
rk1998 n497__vddio n585__vddio 210.6e-3
rk1999 n585__vddio n496__vddio 955.4e-3
rk2000 n496__vddio n586__vddio 557.3e-3
rk2001 n586__vddio n493__vddio 730.7e-3
rk2002 n493__vddio n587__vddio 766e-3
rk2003 n587__vddio n584__vddio 16.4166
rk2004 n551__vddio n588__vddio 692.8e-3
rk2005 n588__vddio n491__vddio 6.215e-3
rk2006 n552__vddio n589__vddio 692.8e-3
rk2007 n589__vddio n485__vddio 6.215e-3
rk2008 n554__vddio n479__vddio 605.7e-3
rk2009 n479__vddio n591__vddio 209e-3
rk2010 n591__vddio n478__vddio 953.9e-3
rk2011 n478__vddio n592__vddio 555.8e-3
rk2012 n592__vddio n475__vddio 729.1e-3
rk2013 n475__vddio n593__vddio 764.4e-3
rk2014 n593__vddio n590__vddio 16.4166
rk2015 n555__vddio n473__vddio 607.3e-3
rk2016 n473__vddio n595__vddio 210.6e-3
rk2017 n595__vddio n472__vddio 955.4e-3
rk2018 n472__vddio n596__vddio 557.3e-3
rk2019 n596__vddio n469__vddio 730.7e-3
rk2020 n469__vddio n597__vddio 766e-3
rk2021 n597__vddio n594__vddio 16.4166
rk2022 n556__vddio n467__vddio 607.3e-3
rk2023 n467__vddio n599__vddio 210.6e-3
rk2024 n599__vddio n466__vddio 955.4e-3
rk2025 n466__vddio n600__vddio 557.3e-3
rk2026 n600__vddio n463__vddio 730.7e-3
rk2027 n463__vddio n601__vddio 766e-3
rk2028 n601__vddio n598__vddio 16.4166
rk2029 n557__vddio n462__vddio 607.4e-3
rk2030 n462__vddio n603__vddio 210.7e-3
rk2031 n603__vddio n459__vddio 955.5e-3
rk2032 n459__vddio n604__vddio 557.4e-3
rk2033 n604__vddio n458__vddio 730.8e-3
rk2034 n458__vddio n605__vddio 766.1e-3
rk2035 n605__vddio n602__vddio 16.4166
rk2036 n559__vddio n456__vddio 607.4e-3
rk2037 n456__vddio n607__vddio 210.7e-3
rk2038 n607__vddio n453__vddio 955.5e-3
rk2039 n453__vddio n608__vddio 557.4e-3
rk2040 n608__vddio n452__vddio 730.8e-3
rk2041 n452__vddio n609__vddio 766.1e-3
rk2042 n609__vddio n606__vddio 16.4166
rk2043 n433__vddio n611__vddio 213.8e-3
rk2044 n611__vddio n432__vddio 958.6e-3
rk2045 n432__vddio n612__vddio 560.6e-3
rk2046 n612__vddio n429__vddio 733.9e-3
rk2047 n429__vddio n613__vddio 769.2e-3
rk2048 n613__vddio n610__vddio 16.4166
rk2049 n588__vddio n615__vddio 296.2e-3
rk2050 n615__vddio n616__vddio 1.041
rk2051 n616__vddio n490__vddio 6.215e-3
rk2052 n589__vddio n618__vddio 296.2e-3
rk2053 n618__vddio n619__vddio 1.041
rk2054 n619__vddio n484__vddio 6.215e-3
rk2055 n616__vddio n620__vddio 642.9e-3
rk2056 n620__vddio n621__vddio 816.3e-3
rk2057 n621__vddio n487__vddio 6.215e-3
rk2058 n619__vddio n622__vddio 642.9e-3
rk2059 n622__vddio n623__vddio 816.3e-3
rk2060 n623__vddio n481__vddio 6.215e-3
rk2061 n621__vddio n624__vddio 851.6e-3
rk2062 n624__vddio n614__vddio 16.4166
rk2063 n623__vddio n625__vddio 851.6e-3
rk2064 n625__vddio n617__vddio 16.4166
rk2065 n535__vddio n536__vddio 3.2632
rk2066 n535__vddio n538__vddio 3.1
rk2067 n535__vddio n540__vddio 3.1
rk2068 n560__vddio n561__vddio 3.1
rk2069 n560__vddio n562__vddio 3.1
rk2070 n560__vddio n563__vddio 3.2632
rk2071 n564__vddio n565__vddio 3.1
rk2072 n564__vddio n566__vddio 3.1
rk2073 n564__vddio n567__vddio 3.2632
rk2074 n568__vddio n569__vddio 3.1
rk2075 n568__vddio n570__vddio 3.1
rk2076 n568__vddio n571__vddio 3.2632
rk2077 n572__vddio n573__vddio 3.1
rk2078 n572__vddio n574__vddio 3.1
rk2079 n572__vddio n575__vddio 3.2632
rk2080 n576__vddio n577__vddio 3.1
rk2081 n576__vddio n578__vddio 3.1
rk2082 n576__vddio n579__vddio 3.2632
rk2083 n580__vddio n581__vddio 3.1
rk2084 n580__vddio n582__vddio 3.1
rk2085 n580__vddio n583__vddio 3.2632
rk2086 n584__vddio n585__vddio 3.1
rk2087 n584__vddio n586__vddio 3.1
rk2088 n584__vddio n587__vddio 3.2632
rk2089 n590__vddio n591__vddio 3.1
rk2090 n590__vddio n592__vddio 3.1
rk2091 n590__vddio n593__vddio 3.2632
rk2092 n594__vddio n595__vddio 3.1
rk2093 n594__vddio n596__vddio 3.1
rk2094 n594__vddio n597__vddio 3.2632
rk2095 n598__vddio n599__vddio 3.1
rk2096 n598__vddio n600__vddio 3.1
rk2097 n598__vddio n601__vddio 3.2632
rk2098 n602__vddio n603__vddio 3.1
rk2099 n602__vddio n604__vddio 3.1
rk2100 n602__vddio n605__vddio 3.2632
rk2101 n606__vddio n607__vddio 3.1
rk2102 n606__vddio n608__vddio 3.1
rk2103 n606__vddio n609__vddio 3.2632
rk2104 n610__vddio n611__vddio 3.1
rk2105 n610__vddio n612__vddio 3.1
rk2106 n610__vddio n613__vddio 3.2632
rk2107 n614__vddio n615__vddio 3.1
rk2108 n617__vddio n618__vddio 3.1
rk2109 n614__vddio n620__vddio 3.1
rk2110 n617__vddio n622__vddio 3.1
rk2111 n614__vddio n624__vddio 3.2632
rk2112 n617__vddio n625__vddio 3.2632
rk2113 n3__i2__net1 n6__i2__net1 1.2339
rk2114 n6__i2__net1 n7__i2__net1 75.5472
rk2115 n5__i2__net1 n6__i2__net1 31
rk2116 n3__i1__net1 n6__i1__net1 1.2339
rk2117 n6__i1__net1 n7__i1__net1 75.5498
rk2118 n5__i1__net1 n6__i1__net1 31
rk2119 n3__i0__net1 n6__i0__net1 1.2339
rk2120 n6__i0__net1 n7__i0__net1 75.5472
rk2121 n5__i0__net1 n6__i0__net1 31
rk2122 n3__i13__i19__i4__net2 n4__i13__i19__i4__net2 75.0403
rk2123 n4__i13__i19__i4__net2 n5__i13__i19__i4__net2 31.3601
rk2124 n3__i13__i18__i4__net2 n4__i13__i18__i4__net2 31.3601
rk2125 n4__i13__i18__i4__net2 n5__i13__i18__i4__net2 75.0403
rk2126 n16__i13__net11 n17__i13__net11 75.4527
rk2127 n17__i13__net11 n18__i13__net11 62.0153
rk2128 n20__i13__net12 n21__i13__net12 75.4527
rk2129 n21__i13__net12 n22__i13__net12 62.0153
rk2130 n10__i13__net1 n21__i13__net1 55.48e-3
rk2131 n21__i13__net1 n19__i13__net1 490.2e-3
rk2132 n10__i13__net2 n25__i13__net2 55.48e-3
rk2133 n25__i13__net2 n23__i13__net2 490.2e-3
rk2134 n6__i13__i19__i4__net2 n2__i13__i19__i4__net2 3.514e-3
rk2135 n2__i13__i18__i4__net2 n6__i13__i18__i4__net2 3.514e-3
rk2136 n11__i13__net18 n13__i13__net18 75.4649
rk2137 n13__i13__net18 n14__i13__net18 519.5e-3
rk2138 n12__i13__net18 n13__i13__net18 62
rk2139 r0 n3__r0 75.4649
rk2140 n3__r0 n4__r0 519.9e-3
rk2141 n2__r0 n3__r0 62
rk2142 n22__i13__net1 n23__i13__net1 31.6782
rk2143 n26__i13__net2 n27__i13__net2 31.6782
rk2144 n7__i13__i19__i4__net2 n8__i13__i19__i4__net2 6.35e-3
rk2145 n9__i13__i19__i4__net2 n11__i13__i19__i4__net2 6.35e-3
rk2146 n8__i13__i19__i4__net2 n9__i13__i19__i4__net2 28.4e-3
rk2147 n10__i13__i19__i4__net2 n11__i13__i19__i4__net2 75
rk2148 n7__i13__i18__i4__net2 n9__i13__i18__i4__net2 6.35e-3
rk2149 n10__i13__i18__i4__net2 n11__i13__i18__i4__net2 6.35e-3
rk2150 n7__i13__i18__i4__net2 n11__i13__i18__i4__net2 28.4e-3
rk2151 n8__i13__i18__i4__net2 n9__i13__i18__i4__net2 75
rk2152 n7__i13__net11 n20__i13__net11 212.1e-3
rk2153 n7__i13__net12 n24__i13__net12 212.1e-3
rk2154 i2__net73 n2__i2__net73 62.4304
rk2155 n2__i2__net73 n3__i2__net73 530.6e-3
rk2156 n3__i2__net73 n4__i2__net73 37.7009
rk2157 n2__i2__net73 n5__i2__net73 75.1559
rk2158 n3__i2__net73 n6__i2__net73 15.7865
rk2159 i1__net73 n2__i1__net73 75.1559
rk2160 n2__i1__net73 n3__i1__net73 530.6e-3
rk2161 n3__i1__net73 n4__i1__net73 15.7865
rk2162 n2__i1__net73 n5__i1__net73 62.4304
rk2163 n3__i1__net73 n6__i1__net73 37.7009
rk2164 i0__net73 n2__i0__net73 62.4304
rk2165 n2__i0__net73 n3__i0__net73 530.6e-3
rk2166 n3__i0__net73 n4__i0__net73 37.7009
rk2167 n2__i0__net73 n5__i0__net73 75.1559
rk2168 n3__i0__net73 n6__i0__net73 15.7865
rk2169 n15__i13__net18 n17__i13__net18 75.3453
rk2170 n17__i13__net18 n18__i13__net18 561.7e-3
rk2171 n16__i13__net18 n17__i13__net18 31
rk2172 n6__r0 n7__r0 561.7e-3
rk2173 n6__r0 n8__r0 75.3453
rk2174 n5__r0 n6__r0 31
rk2175 n2__i18__net3 n31__i18__net3 45.5
rk2176 n38__ck_buff n16__ck_buff 509.5e-3
rk2177 n35__ck_b n19__ck_b 509.5e-3
rk2178 n21__ck_b n36__ck_b 509.5e-3
rk2179 n18__ck_buff n39__ck_buff 509.5e-3
rk2180 n40__ck_buff n20__ck_buff 509.5e-3
rk2181 n37__ck_b n23__ck_b 509.5e-3
rk2182 n152__i18__net4 n153__i18__net4 5.637
rk2183 n153__i18__net4 n154__i18__net4 43.48e-3
rk2185 n152__i18__net4 n153__i18__net4 3.75
rk2186 n156__i18__net4 n157__i18__net4 6.2303
rk2187 n157__i18__net4 n158__i18__net4 177.6e-3
rk2188 n158__i18__net4 n156__i18__net4 4.641
rk2189 n156__i18__net4 n158__i18__net4 3.1
rk2190 n8__i2__net74 n10__i2__net74 75.3852
rk2191 n10__i2__net74 n11__i2__net74 51.22e-3
rk2192 n11__i2__net74 n12__i2__net74 75.4403
rk2193 n11__i2__net74 n13__i2__net74 62.2822
rk2194 n9__i2__net74 n10__i2__net74 62
rk2195 n8__i1__net74 n10__i1__net74 75.3825
rk2196 n10__i1__net74 n11__i1__net74 51.22e-3
rk2197 n11__i1__net74 n12__i1__net74 62.2704
rk2198 n11__i1__net74 n13__i1__net74 75.4286
rk2199 n9__i1__net74 n10__i1__net74 62
rk2200 n8__i0__net74 n10__i0__net74 75.3852
rk2201 n10__i0__net74 n11__i0__net74 51.22e-3
rk2202 n11__i0__net74 n12__i0__net74 75.4403
rk2203 n11__i0__net74 n13__i0__net74 62.2833
rk2204 n9__i0__net74 n10__i0__net74 62
rk2205 n5__i18__net3 n33__i18__net3 45.5
rk2206 i2__net75 n4__i2__net75 45.8942
rk2207 i1__net75 n4__i1__net75 45.8942
rk2208 i0__net75 n4__i0__net75 45.8942
rk2209 n8__i18__net3 n35__i18__net3 45.5
rk2210 n5__i13__i20__net1 n6__i13__i20__net1 31.5319
rk2211 n4__i13__net3 n5__i13__net3 75.5
rk2212 n3__i13__net7 n14__i13__net7 513.2e-3
rk2213 n3__i13__net17 n9__i13__net17 512.4e-3
rk2214 n163__i18__net4 n164__i18__net4 5.637
rk2215 n164__i18__net4 n165__i18__net4 31.89e-3
rk2217 n163__i18__net4 n164__i18__net4 3.75
rk2218 n167__i18__net4 n168__i18__net4 6.2175
rk2219 n168__i18__net4 n169__i18__net4 190.5e-3
rk2220 n169__i18__net4 n167__i18__net4 4.641
rk2221 n167__i18__net4 n169__i18__net4 3.1
rk2222 n41__ck_buff n42__ck_buff 1.213
rk2223 n43__ck_buff n44__ck_buff 1.213
rk2224 n45__ck_buff n46__ck_buff 1.213
rk2225 n11__i18__net3 n36__i18__net3 45.5
rk2226 n3__i13__net23 n5__i13__net23 512.1e-3
rk2227 n3__i13__net18 n20__i13__net18 511.3e-3
rk2228 n41__ck_b n38__ck_b 1.2288
rk2229 n42__ck_b n39__ck_b 1.2288
rk2230 n43__ck_b n40__ck_b 1.2288
rk2231 n14__i2__net74 n15__i2__net74 75.812
rk2232 n14__i1__net74 n15__i1__net74 75.812
rk2233 n14__i0__net74 n15__i0__net74 75.812
rk2234 n14__i18__net3 n39__i18__net3 45
rk2235 n30__reset_buff n33__reset_buff 4.237e-3
rk2236 n34__reset_buff n20__reset_buff 4.237e-3
rk2237 n33__reset_buff n34__reset_buff 23.66e-3
rk2238 n35__reset_buff n22__reset_buff 4.237e-3
rk2239 n31__reset_buff n36__reset_buff 4.237e-3
rk2240 n35__reset_buff n36__reset_buff 23.66e-3
rk2241 n32__reset_buff n37__reset_buff 4.237e-3
rk2242 n38__reset_buff n24__reset_buff 4.237e-3
rk2243 n37__reset_buff n38__reset_buff 23.66e-3
rk2244 n8__i13__i20__net1 n9__i13__i20__net1 37.7009
rk2245 n9__i13__i20__net1 n7__i13__i20__net1 283.1e-3
rk2246 n7__i13__i20__net1 n10__i13__i20__net1 31
rk2247 n9__i13__i20__net1 n3__i13__i20__net1 170.8e-3
rk2248 n7__i13__net3 n8__i13__net3 15.7843
rk2249 n8__i13__net3 n6__i13__net3 238.6e-3
rk2250 n6__i13__net3 n9__i13__net3 75
rk2251 n8__i13__net3 n2__i13__net3 45.1981
rk2252 n180__i18__net4 n181__i18__net4 5.637
rk2253 n181__i18__net4 n178__i18__net4 40.59e-3
rk2255 n180__i18__net4 n181__i18__net4 3.75
rk2256 n183__i18__net4 n179__i18__net4 6.2271
rk2257 n179__i18__net4 n184__i18__net4 180.8e-3
rk2258 n184__i18__net4 n183__i18__net4 4.641
rk2259 n183__i18__net4 n184__i18__net4 3.1
rk2260 n6__i13__net23 n8__i13__net23 554.6e-3
rk2261 n8__i13__net23 n9__i13__net23 31.3424
rk2262 n7__i13__net23 n8__i13__net23 75
rk2263 r2 n2__r2 31.1559
rk2264 n2__r2 n3__r2 75.1687
rk2265 n17__i18__net3 n41__i18__net3 45.5
rk2266 n4__i2__net74 n16__i2__net74 228.1e-3
rk2267 n4__i1__net74 n16__i1__net74 228.1e-3
rk2268 n4__i0__net74 n16__i0__net74 228.1e-3
rk2269 n20__i18__net3 n43__i18__net3 45.5
rk2270 n7__i13__net18 n22__i13__net18 6.854e-3
rk2271 n185__i18__net4 n186__i18__net4 5.637
rk2272 n186__i18__net4 n187__i18__net4 43.48e-3
rk2274 n185__i18__net4 n186__i18__net4 3.75
rk2275 n189__i18__net4 n190__i18__net4 6.2303
rk2276 n190__i18__net4 n191__i18__net4 177.6e-3
rk2277 n191__i18__net4 n189__i18__net4 4.641
rk2278 n189__i18__net4 n191__i18__net4 3.1
rk2279 n3__i13__i20__i4__net2 n4__i13__i20__i4__net2 75.0403
rk2280 n4__i13__i20__i4__net2 n5__i13__i20__i4__net2 31.3601
rk2281 n6__i2__net75 n7__i2__net75 62.4304
rk2282 n7__i2__net75 n8__i2__net75 277e-3
rk2283 n8__i2__net75 n9__i2__net75 37.7116
rk2284 n7__i2__net75 n10__i2__net75 75.1559
rk2285 n8__i2__net75 n12__i2__net75 307.9e-3
rk2286 n12__i2__net75 n5__i2__net75 112.8e-3
rk2287 n11__i2__net75 n12__i2__net75 15.5
rk2288 n6__i1__net75 n7__i1__net75 75.1559
rk2289 n7__i1__net75 n8__i1__net75 277e-3
rk2290 n8__i1__net75 n10__i1__net75 307.9e-3
rk2291 n7__i1__net75 n11__i1__net75 62.4304
rk2292 n8__i1__net75 n12__i1__net75 37.7116
rk2293 n10__i1__net75 n5__i1__net75 108e-3
rk2294 n9__i1__net75 n10__i1__net75 15.5
rk2295 n6__i0__net75 n7__i0__net75 62.4304
rk2296 n7__i0__net75 n8__i0__net75 277e-3
rk2297 n8__i0__net75 n9__i0__net75 37.7116
rk2298 n7__i0__net75 n10__i0__net75 75.1559
rk2299 n8__i0__net75 n12__i0__net75 307.9e-3
rk2300 n12__i0__net75 n5__i0__net75 112.8e-3
rk2301 n11__i0__net75 n12__i0__net75 15.5
rk2302 n23__i18__net3 n45__i18__net3 45.5
rk2303 n16__i13__net7 n17__i13__net7 75.4527
rk2304 n17__i13__net7 n18__i13__net7 62.0153
rk2305 n10__i13__net18 n23__i13__net18 55.48e-3
rk2306 n23__i13__net18 n24__i13__net18 990.2e-3
rk2307 n6__i13__i20__i4__net2 n2__i13__i20__i4__net2 3.514e-3
rk2308 n44__ck_b n25__ck_b 509.5e-3
rk2309 n47__ck_buff n28__ck_buff 509.5e-3
rk2310 n30__ck_buff n48__ck_buff 509.5e-3
rk2311 n27__ck_b n45__ck_b 509.5e-3
rk2312 n46__ck_b n29__ck_b 509.5e-3
rk2313 n49__ck_buff n32__ck_buff 509.5e-3
rk2314 n5__r1 n7__r1 75.4649
rk2315 n7__r1 n8__r1 519.5e-3
rk2316 n6__r1 n7__r1 62
rk2317 n26__i18__net3 n46__i18__net3 45.5
rk2318 n8__i2__net76 n10__i2__net76 75.3852
rk2319 n10__i2__net76 n11__i2__net76 51.22e-3
rk2320 n11__i2__net76 n12__i2__net76 75.4403
rk2321 n11__i2__net76 n13__i2__net76 62.2822
rk2322 n9__i2__net76 n10__i2__net76 62
rk2323 n8__i1__net76 n10__i1__net76 75.3825
rk2324 n10__i1__net76 n11__i1__net76 51.22e-3
rk2325 n11__i1__net76 n12__i1__net76 62.2704
rk2326 n11__i1__net76 n13__i1__net76 75.4286
rk2327 n9__i1__net76 n10__i1__net76 62
rk2328 n8__i0__net76 n10__i0__net76 75.3852
rk2329 n10__i0__net76 n11__i0__net76 51.22e-3
rk2330 n11__i0__net76 n12__i0__net76 75.4403
rk2331 n11__i0__net76 n13__i0__net76 62.2833
rk2332 n9__i0__net76 n10__i0__net76 62
rk2333 n196__i18__net4 n197__i18__net4 5.637
rk2334 n197__i18__net4 n198__i18__net4 31.89e-3
rk2336 n196__i18__net4 n197__i18__net4 3.75
rk2337 n200__i18__net4 n201__i18__net4 6.2175
rk2338 n201__i18__net4 n202__i18__net4 190.5e-3
rk2339 n202__i18__net4 n200__i18__net4 4.641
rk2340 n200__i18__net4 n202__i18__net4 3.1
rk2341 n26__i13__net18 n27__i13__net18 31.6782
rk2342 n7__i13__i20__i4__net2 n8__i13__i20__i4__net2 6.35e-3
rk2343 n9__i13__i20__i4__net2 n11__i13__i20__i4__net2 6.35e-3
rk2344 n8__i13__i20__i4__net2 n9__i13__i20__i4__net2 28.4e-3
rk2345 n10__i13__i20__i4__net2 n11__i13__i20__i4__net2 75
rk2346 n7__i13__net7 n20__i13__net7 212.1e-3
rk2347 i2__net77 n7__i2__net77 45.8942
rk2348 i1__net77 n7__i1__net77 45.8942
rk2349 i0__net77 n7__i0__net77 45.8942
rk2350 n9__r1 n11__r1 75.3453
rk2351 n11__r1 n12__r1 561.7e-3
rk2352 n10__r1 n11__r1 31
rk2355 n624__vss n625__vss 1.0383
rk2356 n625__vss n626__vss 174.4e-3
rk2357 n626__vss n627__vss 329.9e-3
rk2358 n627__vss n628__vss 354.2e-3
rk2359 n624__vss n623__vss 5.2204
rk2360 n626__vss n630__vss 887.9e-3
rk2361 n630__vss n629__vss 5.2204
rk2362 n627__vss n632__vss 887.9e-3
rk2363 n632__vss n631__vss 5.2204
rk2364 n628__vss n634__vss 898.9e-3
rk2365 n634__vss n633__vss 5.2204
rk2366 n628__vss n635__vss 306.9e-3
rk2367 n635__vss n637__vss 887.9e-3
rk2368 n637__vss n636__vss 5.2204
rk2369 n635__vss n639__vss 1.2193
rk2370 n639__vss n638__vss 5.2204
rk2371 n623__vss n624__vss 4.1667
rk2372 n629__vss n630__vss 4.1667
rk2373 n631__vss n632__vss 4.1667
rk2374 n633__vss n634__vss 4.1667
rk2375 n636__vss n637__vss 4.1667
rk2376 n638__vss n639__vss 4.1667
rk2377 n636__vddio n637__vddio 6.4123
rk2378 n637__vddio n638__vddio 1.541
rk2379 n638__vddio n639__vddio 1.2085
rk2380 n639__vddio n640__vddio 174.4e-3
rk2381 n640__vddio n641__vddio 329.9e-3
rk2382 n641__vddio n642__vddio 354.2e-3
rk2383 n640__vddio n644__vddio 1.058
rk2384 n644__vddio n645__vddio 1.541
rk2385 n645__vddio n643__vddio 6.4123
rk2386 n641__vddio n647__vddio 1.058
rk2387 n647__vddio n648__vddio 1.541
rk2388 n648__vddio n646__vddio 6.4123
rk2389 n642__vddio n649__vddio 306.9e-3
rk2390 n649__vddio n651__vddio 1.3894
rk2391 n651__vddio n652__vddio 1.541
rk2392 n652__vddio n650__vddio 6.4123
rk2393 n642__vddio n654__vddio 1.0691
rk2394 n654__vddio n655__vddio 1.541
rk2395 n655__vddio n653__vddio 6.4123
rk2396 n649__vddio n657__vddio 1.058
rk2397 n657__vddio n658__vddio 1.541
rk2398 n658__vddio n656__vddio 6.4123
rk2399 n636__vddio n637__vddio 3.1
rk2400 n636__vddio n638__vddio 3.1
rk2401 n643__vddio n644__vddio 3.1
rk2402 n643__vddio n645__vddio 3.1
rk2403 n646__vddio n647__vddio 3.1
rk2404 n646__vddio n648__vddio 3.1
rk2405 n650__vddio n651__vddio 3.1
rk2406 n650__vddio n652__vddio 3.1
rk2407 n653__vddio n654__vddio 3.1
rk2408 n653__vddio n655__vddio 3.1
rk2409 n656__vddio n657__vddio 3.1
rk2410 n656__vddio n658__vddio 3.1
rk2411 n16__reset_b n25__reset_b 40.14e-3
rk2412 n18__reset_b n26__reset_b 40.14e-3
rk2413 n20__reset_b n27__reset_b 40.14e-3
rk2416 n640__vss n641__vss 4.9167
rk2417 n641__vss n642__vss 574.2e-3
rk2418 n642__vss n643__vss 574.2e-3
rk2419 n643__vss n644__vss 93.1e-3
rk2420 n644__vss n645__vss 97.67e-3
rk2421 n645__vss n646__vss 133.6e-3
rk2422 n646__vss n647__vss 248.6e-3
rk2423 n647__vss n648__vss 219.9e-3
rk2424 n648__vss n649__vss 194.6e-3
rk2425 n649__vss n650__vss 33.28e-3
rk2426 n650__vss n651__vss 64.39e-3
rk2427 n651__vss n652__vss 139.5e-3
rk2428 n652__vss n653__vss 33.28e-3
rk2429 n653__vss n654__vss 64.39e-3
rk2430 n654__vss n655__vss 159.9e-3
rk2431 n655__vss n656__vss 97.67e-3
rk2432 n656__vss n657__vss 97.88e-3
rk2433 n657__vss n658__vss 97.88e-3
rk2434 n658__vss n659__vss 110.8e-3
rk2435 n659__vss n660__vss 132.4e-3
rk2436 n660__vss n661__vss 145.7e-3
rk2437 n644__vss n662__vss 37.6834
rk2438 n645__vss n663__vss 37.6727
rk2439 n646__vss n664__vss 75.207
rk2440 n648__vss n665__vss 75.207
rk2441 n649__vss n666__vss 75.207
rk2442 n651__vss n667__vss 75.2123
rk2443 n652__vss n668__vss 37.6727
rk2444 n654__vss n669__vss 37.6834
rk2445 n655__vss n670__vss 37.6727
rk2446 n656__vss n671__vss 37.6834
rk2447 n657__vss n672__vss 37.6798
rk2448 n658__vss n673__vss 37.6727
rk2449 n659__vss n674__vss 37.6727
rk2450 n660__vss n675__vss 37.6829
rk2451 n661__vss n676__vss 37.6691
rk2452 n661__vss n677__vss 88.31e-3
rk2453 n677__vss n678__vss 37.6834
rk2454 n677__vss n402__vss 51.23e-3
rk2455 n402__vss n679__vss 37.6798
rk2456 n402__vss n680__vss 144.5e-3
rk2457 n680__vss n681__vss 37.6749
rk2458 n680__vss n682__vss 110.8e-3
rk2459 n682__vss n683__vss 37.6727
rk2460 n682__vss n684__vss 110.8e-3
rk2461 n684__vss n685__vss 37.6727
rk2462 n684__vss n686__vss 66.78e-3
rk2463 n686__vss n687__vss 53.62e-3
rk2464 n687__vss n688__vss 37.6727
rk2465 n687__vss n689__vss 110.8e-3
rk2466 n689__vss n690__vss 37.6727
rk2467 n689__vss n691__vss 61.78e-3
rk2468 n691__vss n692__vss 37.6727
rk2469 n691__vss n693__vss 97.67e-3
rk2470 n693__vss n694__vss 37.6727
rk2471 n693__vss n695__vss 79.72e-3
rk2472 n695__vss n696__vss 75.2027
rk2473 n695__vss n697__vss 168.5e-3
rk2474 n697__vss n698__vss 179.2e-3
rk2475 n698__vss n699__vss 37.6727
rk2476 n698__vss n700__vss 97.67e-3
rk2477 n700__vss n701__vss 37.6727
rk2478 n700__vss n702__vss 61.78e-3
rk2479 n702__vss n703__vss 75.207
rk2480 n702__vss n704__vss 110.8e-3
rk2481 n704__vss n705__vss 75.2047
rk2482 n704__vss n706__vss 123e-3
rk2483 n706__vss n707__vss 75.3975
rk2484 n640__vss n641__vss 3.1
rk2485 n640__vss n642__vss 3.1
rk2486 n640__vss n643__vss 3.1
rk2487 n640__vss n647__vss 3.1
rk2488 n640__vss n650__vss 20.6667
rk2489 n640__vss n653__vss 20.6667
rk2490 n640__vss n657__vss 4.4286
rk2491 n640__vss n661__vss 3.1
rk2492 n640__vss n686__vss 3.1
rk2493 n640__vss n697__vss 3.1
rk2494 n640__vss n706__vss 3.1
rk2495 n4__i2__net76 n14__i2__net76 212e-3
rk2496 n14__i2__net76 n15__i2__net76 62.0166
rk2497 n4__i1__net76 n14__i1__net76 212e-3
rk2498 n14__i1__net76 n15__i1__net76 62.0166
rk2499 n4__i0__net76 n14__i0__net76 212e-3
rk2500 n14__i0__net76 n15__i0__net76 62.0166
rk2503 n8__i2__net77 n9__i2__net77 37.6937
rk2504 n9__i2__net77 n11__i2__net77 290e-3
rk2505 n11__i2__net77 n12__i2__net77 612.8e-3
rk2506 n10__i2__net77 n11__i2__net77 15.5
rk2507 n8__i1__net77 n9__i1__net77 37.6937
rk2508 n9__i1__net77 n11__i1__net77 290e-3
rk2509 n11__i1__net77 n12__i1__net77 608e-3
rk2510 n10__i1__net77 n11__i1__net77 15.5
rk2511 n8__i0__net77 n9__i0__net77 37.6937
rk2512 n9__i0__net77 n11__i0__net77 290e-3
rk2513 n11__i0__net77 n12__i0__net77 612.8e-3
rk2514 n10__i0__net77 n11__i0__net77 15.5
rk2515 n6__serial_out_b_high n7__serial_out_b_high 31.5698
rk2516 n5__i2__net77 n13__i2__net77 45.5268
rk2517 n5__i1__net77 n13__i1__net77 45.5268
rk2518 n5__i0__net77 n13__i0__net77 45.5268
rk2519 n3__i12__bio n4__i12__bio 38.1033
rk2522 n8__serial_out_b_high n9__serial_out_b_high 37.9387
rk2523 n9__serial_out_b_high n10__serial_out_b_high 38.3822
rk2524 n9__serial_out_b_high n11__serial_out_b_high 1.2679
rk2525 n9__serial_out n20__serial_out 119.8e-3
rk2526 n20__serial_out n21__serial_out 37.708
rk2527 n20__serial_out n22__serial_out 177e-3
rk2528 n22__serial_out n23__serial_out 15.5974
rk2529 n10__net4 n12__net4 119.8e-3
rk2530 n12__net4 n13__net4 177e-3
rk2531 n13__net4 n14__net4 15.5974
rk2532 n12__net4 n15__net4 37.708
rk2533 n8__net3 n10__net3 119.8e-3
rk2534 n10__net3 n11__net3 37.708
rk2535 n10__net3 n12__net3 177e-3
rk2536 n12__net3 n13__net3 15.5974
rk2537 n51__i18__net3 n52__i18__net3 13.5161
rk2538 n52__i18__net3 n53__i18__net3 953.9e-3
rk2539 n53__i18__net3 n54__i18__net3 326.3e-3
rk2540 n54__i18__net3 n49__i18__net3 624e-3
rk2542 n53__i18__net3 n57__i18__net3 831.9e-3
rk2543 n57__i18__net3 n56__i18__net3 4.4901
rk2544 n54__i18__net3 n59__i18__net3 828.3e-3
rk2545 n59__i18__net3 n58__i18__net3 4.4901
rk2546 n54__i18__net3 n61__i18__net3 950.3e-3
rk2547 n61__i18__net3 n60__i18__net3 13.5161
rk2548 n51__i18__net3 n52__i18__net3 3.75
rk2549 n29__i18__net3 n49__i18__net3 45
rk2550 n56__i18__net3 n57__i18__net3 3.875
rk2551 n58__i18__net3 n59__i18__net3 3.875
rk2552 n60__i18__net3 n61__i18__net3 3.75
rk2555 i2__q n2__i2__q 15.8098
rk2556 n2__i2__q n3__i2__q 37.655
rk2557 i1__q n2__i1__q 37.655
rk2558 n2__i1__q n3__i1__q 15.8098
rk2559 i0__q n2__i0__q 15.8098
rk2560 n2__i0__q n3__i0__q 37.655
rk2561 n5__i12__bio n6__i12__bio 31.2929
rk2562 n6__i12__bio n7__i12__bio 518.8e-3
rk2563 n7__i12__bio i12__bio 19.3e-3
rk2564 n6__i12__bio n8__i12__bio 411e-3
rk2565 n8__i12__bio n9__i12__bio 37.6055
rk2566 n709__vss n710__vss 706.6e-3
rk2567 n709__vss n708__vss 4.7661
rk2568 n710__vss n712__vss 393.3e-3
rk2569 n712__vss n711__vss 4.7661
rk2570 n710__vss n714__vss 710.5e-3
rk2571 n714__vss n713__vss 4.7661
rk2572 n708__vss n709__vss 12.5
rk2573 n711__vss n712__vss 12.5
rk2574 n713__vss n714__vss 12.5
rk2575 n659__vddio n660__vddio 5.2651
rk2576 n660__vddio n661__vddio 1.4338
rk2577 n661__vddio n663__vddio 1.4377
rk2578 n663__vddio n662__vddio 5.2651
rk2579 n661__vddio n665__vddio 1.1204
rk2580 n665__vddio n664__vddio 5.2651
rk2581 n659__vddio n660__vddio 3.1
rk2582 n662__vddio n663__vddio 3.1
rk2583 n664__vddio n665__vddio 3.1
rk2584 n12__serial_out_b_high serial_out_b_high 529.6e-3
rk2585 n13__i18__net2 n14__i18__net2 6.0896
rk2586 n14__i18__net2 n2__i18__net2 23.0225
rk2587 n14__i18__net2 n15__i18__net2 4.2396
rk2588 n11__i12__bcore_bar n12__i12__bcore_bar 75.2373
rk2589 n12__i12__bcore_bar n5__i12__bcore_bar 754.7e-3
rk2591 n12__i12__bcore_bar n14__i12__bcore_bar 31.3015
rk2593 n12__r0 n14__r0 570.8e-3
rk2594 n7__r2 n9__r2 556.1e-3
rk2595 n3__r1 n13__r1 573.2e-3
rk2596 n24__serial_out n12__serial_out 23.0098
rk2597 n31__vdd n33__vdd 1.0487
rk2598 n33__vdd n34__vdd 191.2e-3
rk2599 n34__vdd n35__vdd 126.2e-3
rk2600 n35__vdd n36__vdd 110.6e-3
rk2601 n36__vdd n37__vdd 48.62e-3
rk2602 n37__vdd n38__vdd 66.78e-3
rk2603 n38__vdd n39__vdd 449.4e-3
rk2604 n39__vdd n23__vdd 97.49e-3
rk2605 n23__vdd n40__vdd 17.12e-3
rk2606 n40__vdd n41__vdd 109.8e-3
rk2607 n41__vdd n42__vdd 460.2e-3
rk2608 n42__vdd n43__vdd 104.8e-3
rk2609 n43__vdd n44__vdd 126e-3
rk2610 n44__vdd n45__vdd 110.4e-3
rk2611 n45__vdd n46__vdd 230.5e-3
rk2612 n46__vdd n47__vdd 334.5e-3
rk2613 n47__vdd n48__vdd 238.8e-3
rk2614 n48__vdd n49__vdd 277.1e-3
rk2615 n49__vdd n50__vdd 148.7e-3
rk2616 n50__vdd n51__vdd 110.4e-3
rk2617 n51__vdd n52__vdd 35.46e-3
rk2618 n52__vdd n53__vdd 25.89e-3
rk2619 n53__vdd n54__vdd 97.25e-3
rk2620 n54__vdd n55__vdd 110.4e-3
rk2621 n55__vdd n56__vdd 61.36e-3
rk2622 n56__vdd n57__vdd 189.8e-3
rk2623 n57__vdd n58__vdd 64.18e-3
rk2624 n58__vdd n59__vdd 97.25e-3
rk2625 n59__vdd n60__vdd 265.9e-3
rk2626 n60__vdd n61__vdd 144.3e-3
rk2627 n61__vdd n62__vdd 168.3e-3
rk2628 n62__vdd n63__vdd 110.4e-3
rk2629 n63__vdd n64__vdd 61.36e-3
rk2630 n64__vdd n65__vdd 97.25e-3
rk2631 n65__vdd n66__vdd 110.4e-3
rk2632 n66__vdd n67__vdd 22.3e-3
rk2633 n67__vdd n5__vdd 82.54e-3
rk2634 n34__vdd n68__vdd 31.3268
rk2635 n35__vdd n69__vdd 31.4136
rk2636 n35__vdd n70__vdd 31.4136
rk2637 n36__vdd n71__vdd 31.1841
rk2638 n37__vdd n72__vdd 15.7583
rk2639 n39__vdd n73__vdd 31.4136
rk2640 n39__vdd n74__vdd 31.4136
rk2641 n40__vdd n75__vdd 31.3078
rk2642 n40__vdd n76__vdd 31.3078
rk2643 n41__vdd n77__vdd 31.2709
rk2644 n41__vdd n78__vdd 31.2709
rk2645 n43__vdd n79__vdd 31.4136
rk2646 n43__vdd n80__vdd 31.4136
rk2647 n44__vdd n81__vdd 31.4136
rk2648 n44__vdd n82__vdd 31.4136
rk2649 n45__vdd n83__vdd 31.2709
rk2650 n45__vdd n84__vdd 31.2709
rk2651 n47__vdd n85__vdd 31.4136
rk2652 n47__vdd n86__vdd 31.4136
rk2653 n49__vdd n87__vdd 31.4136
rk2654 n49__vdd n88__vdd 31.4136
rk2655 n50__vdd n89__vdd 15.8451
rk2656 n50__vdd n90__vdd 15.8451
rk2657 n51__vdd n91__vdd 15.8451
rk2658 n51__vdd n92__vdd 15.8451
rk2659 n53__vdd n93__vdd 15.8451
rk2660 n53__vdd n94__vdd 15.8451
rk2661 n54__vdd n95__vdd 15.8451
rk2662 n54__vdd n96__vdd 15.8451
rk2663 n55__vdd n97__vdd 62.4486
rk2664 n55__vdd n98__vdd 62.4486
rk2665 n56__vdd n99__vdd 62.4771
rk2666 n56__vdd n100__vdd 62.4771
rk2667 n58__vdd n101__vdd 15.8451
rk2668 n58__vdd n102__vdd 15.8451
rk2669 n59__vdd n103__vdd 15.8451
rk2670 n59__vdd n104__vdd 15.8451
rk2671 n60__vdd n105__vdd 62.5087
rk2672 n60__vdd n106__vdd 62.5087
rk2673 n62__vdd n107__vdd 15.8451
rk2674 n62__vdd n108__vdd 15.8451
rk2675 n63__vdd n109__vdd 15.8451
rk2676 n63__vdd n110__vdd 15.8451
rk2677 n64__vdd n111__vdd 15.8451
rk2678 n64__vdd n112__vdd 15.8451
rk2679 n65__vdd n113__vdd 15.8451
rk2680 n65__vdd n114__vdd 15.8451
rk2681 n66__vdd n115__vdd 62.4486
rk2682 n66__vdd n116__vdd 62.4486
rk2683 n5__vdd n117__vdd 62.3867
rk2684 n5__vdd n118__vdd 211.3e-3
rk2685 n118__vdd n119__vdd 15.8451
rk2686 n5__vdd n120__vdd 62.3867
rk2687 n118__vdd n121__vdd 97.25e-3
rk2688 n121__vdd n122__vdd 15.8451
rk2689 n118__vdd n123__vdd 15.8451
rk2690 n121__vdd n124__vdd 181.4e-3
rk2691 n124__vdd n125__vdd 84.51e-3
rk2692 n125__vdd n126__vdd 62.5087
rk2693 n121__vdd n127__vdd 15.8451
rk2695 n125__vdd n129__vdd 62.5087
rk2696 n32__vdd n33__vdd 4.1667
rk2697 n32__vdd n38__vdd 3.75
rk2698 n32__vdd n40__vdd 3.75
rk2699 n32__vdd n42__vdd 3.75
rk2700 n32__vdd n46__vdd 3.75
rk2701 n32__vdd n48__vdd 3.75
rk2702 n32__vdd n52__vdd 5.3571
rk2703 n32__vdd n57__vdd 3.75
rk2704 n32__vdd n61__vdd 3.75
rk2705 n32__vdd n67__vdd 3.75
rk2706 n32__vdd n124__vdd 3.75
rk2707 n130__vdd n131__vdd 31.2204
rk2708 n131__vdd n132__vdd 25.0014
rk2709 n5__net7 n11__net7 176e-3
rk2710 n11__net7 n12__net7 75.1652
rk2711 n11__net7 n13__net7 31.208
rk2712 n5__net6 n11__net6 176e-3
rk2713 n11__net6 n12__net6 31.208
rk2714 n11__net6 n13__net6 75.1652
rk2715 n5__net8 n11__net8 176e-3
rk2716 n11__net8 n12__net8 75.1652
rk2717 n11__net8 n13__net8 31.208
rk2718 n670__vddio n671__vddio 504.2e-3
rk2719 n671__vddio n673__vddio 21.32e-3
rk2720 n673__vddio n674__vddio 241.4e-3
rk2722 n671__vddio n676__vddio 31.3632
rk2723 n674__vddio n677__vddio 31.3632
rk2724 n672__vddio n673__vddio 25
rk2725 n13__serial_out_b_high n3__serial_out_b_high 11.8517
rk2726 n7__i18__net1 n8__i18__net1 9.857
rk2727 n8__i18__net1 n2__i18__net1 23.0933
rk2728 n8__i18__net1 n9__i18__net1 6.2725
rk2729 n8__r0_buff n9__r0_buff 31.209
rk2730 n9__r0_buff n10__r0_buff 171.3e-3
rk2731 n10__r0_buff n11__r0_buff 75.1706
rk2732 n9__r0_buff n12__r0_buff 89.05e-3
rk2733 n12__r0_buff n13__r0_buff 75.0754
rk2734 n10__r0_buff n14__r0_buff 31.2187
rk2735 n8__r2_buff n9__r2_buff 31.1838
rk2736 n9__r2_buff n10__r2_buff 104.5e-3
rk2737 n10__r2_buff n12__r2_buff 37.69e-3
rk2738 n9__r2_buff n13__r2_buff 171.3e-3
rk2739 n13__r2_buff n14__r2_buff 31.2187
rk2740 n13__r2_buff n15__r2_buff 75.1706
rk2741 n11__r2_buff n12__r2_buff 75
rk2742 n8__r1_buff n9__r1_buff 31.209
rk2743 n9__r1_buff n10__r1_buff 171.3e-3
rk2744 n10__r1_buff n11__r1_buff 75.1706
rk2745 n9__r1_buff n12__r1_buff 89.05e-3
rk2746 n12__r1_buff n13__r1_buff 75.0754
rk2747 n10__r1_buff n14__r1_buff 31.2187
rk2748 n133__vdd n135__vdd 31.4088
rk2749 n135__vdd n136__vdd 33.28e-3
rk2750 n136__vdd n137__vdd 107.5e-3
rk2751 n137__vdd n138__vdd 23.71e-3
rk2752 n138__vdd n139__vdd 404.7e-3
rk2753 n139__vdd n140__vdd 27.62e-3
rk2754 n140__vdd n141__vdd 75.46e-3
rk2755 n141__vdd n142__vdd 57.47e-3
rk2756 n142__vdd n143__vdd 90.84e-3
rk2757 n143__vdd n144__vdd 103.1e-3
rk2758 n144__vdd n145__vdd 18.72e-3
rk2759 n145__vdd n146__vdd 38.75e-3
rk2760 n146__vdd n147__vdd 236.6e-3
rk2761 n147__vdd n148__vdd 90.84e-3
rk2762 n148__vdd n149__vdd 166.7e-3
rk2763 n149__vdd n150__vdd 81.02e-3
rk2764 n150__vdd n151__vdd 419e-3
rk2765 n151__vdd n152__vdd 1.0449
rk2766 n152__vdd n153__vdd 120.2e-3
rk2767 n153__vdd n154__vdd 97.67e-3
rk2768 n154__vdd n155__vdd 61.99e-3
rk2769 n155__vdd n156__vdd 35.68e-3
rk2770 n156__vdd n157__vdd 149.1e-3
rk2771 n157__vdd n158__vdd 27.09e-3
rk2772 n158__vdd n159__vdd 50.03e-3
rk2773 n159__vdd n160__vdd 33.28e-3
rk2774 n160__vdd n161__vdd 13.93e-3
rk2775 n161__vdd n162__vdd 47.42e-3
rk2776 n162__vdd n163__vdd 84.57e-3
rk2777 n163__vdd n164__vdd 14.05e-3
rk2778 n164__vdd n165__vdd 109.7e-3
rk2779 n165__vdd n166__vdd 61.78e-3
rk2780 n166__vdd n167__vdd 63.19e-3
rk2781 n167__vdd n168__vdd 191.2e-3
rk2782 n168__vdd n169__vdd 28.28e-3
rk2783 n169__vdd n170__vdd 68.96e-3
rk2784 n170__vdd n171__vdd 125.2e-3
rk2785 n171__vdd n172__vdd 33.28e-3
rk2786 n172__vdd n173__vdd 64.39e-3
rk2787 n173__vdd n174__vdd 42.64e-3
rk2788 n174__vdd n175__vdd 96.47e-3
rk2789 n175__vdd n176__vdd 47.64e-3
rk2790 n176__vdd n177__vdd 50.03e-3
rk2791 n177__vdd n178__vdd 159.7e-3
rk2792 n178__vdd n179__vdd 97.25e-3
rk2793 n179__vdd n180__vdd 97.67e-3
rk2794 n180__vdd n181__vdd 97.67e-3
rk2795 n181__vdd n182__vdd 56.78e-3
rk2796 n182__vdd n183__vdd 53.41e-3
rk2797 n183__vdd n184__vdd 43.84e-3
rk2798 n184__vdd n185__vdd 85.82e-3
rk2799 n185__vdd n186__vdd 14.15e-3
rk2800 n186__vdd n187__vdd 95.39e-3
rk2801 n187__vdd n188__vdd 38.07e-3
rk2802 n188__vdd n189__vdd 88.31e-3
rk2803 n189__vdd n190__vdd 35.46e-3
rk2804 n190__vdd n191__vdd 61.57e-3
rk2805 n191__vdd n192__vdd 97.46e-3
rk2806 n192__vdd n193__vdd 61.78e-3
rk2807 n193__vdd n194__vdd 48.05e-3
rk2808 n194__vdd n195__vdd 13.99e-3
rk2809 n195__vdd n196__vdd 97.1e-3
rk2810 n196__vdd n197__vdd 66.78e-3
rk2811 n197__vdd n198__vdd 53.41e-3
rk2812 n198__vdd n199__vdd 110.4e-3
rk2813 n199__vdd n200__vdd 61.36e-3
rk2814 n200__vdd n201__vdd 97.25e-3
rk2815 n201__vdd n202__vdd 110.4e-3
rk2816 n202__vdd n203__vdd 61.36e-3
rk2817 n203__vdd n204__vdd 74.94e-3
rk2818 n204__vdd n1__vdd 82.54e-3
rk2819 n1__vdd n205__vdd 96.48e-3
rk2820 n205__vdd n206__vdd 97.25e-3
rk2821 n206__vdd n207__vdd 265.9e-3
rk2822 n207__vdd n208__vdd 29.48e-3
rk2823 n208__vdd n209__vdd 266.9e-3
rk2824 n209__vdd n210__vdd 31.2111
rk2825 n136__vdd n211__vdd 31.3268
rk2826 n138__vdd n212__vdd 31.3268
rk2827 n139__vdd n213__vdd 15.7599
rk2828 n141__vdd n214__vdd 15.7599
rk2829 n142__vdd n215__vdd 15.7599
rk2830 n143__vdd n216__vdd 15.7599
rk2831 n144__vdd n217__vdd 62.3633
rk2832 n146__vdd n218__vdd 62.3919
rk2833 n147__vdd n219__vdd 15.7599
rk2834 n148__vdd n220__vdd 15.7599
rk2835 n150__vdd n221__vdd 62.4263
rk2836 n151__vdd n222__vdd 15.7599
rk2837 n152__vdd n223__vdd 31.191
rk2838 n153__vdd n224__vdd 20.8822
rk2839 n154__vdd n225__vdd 20.8982
rk2840 n156__vdd n226__vdd 20.8822
rk2841 n157__vdd n227__vdd 15.7583
rk2842 n158__vdd n228__vdd 15.7797
rk2843 n160__vdd n229__vdd 15.7583
rk2844 n161__vdd n230__vdd 15.7583
rk2845 n162__vdd n231__vdd 15.7583
rk2846 n163__vdd n232__vdd 31.3317
rk2847 n164__vdd n233__vdd 15.761
rk2848 n165__vdd n234__vdd 62.3618
rk2849 n166__vdd n235__vdd 62.3903
rk2850 n168__vdd n236__vdd 15.7583
rk2851 n169__vdd n237__vdd 31.3268
rk2852 n170__vdd n238__vdd 15.7583
rk2853 n171__vdd n239__vdd 31.3268
rk2854 n173__vdd n240__vdd 31.3375
rk2855 n174__vdd n241__vdd 62.4219
rk2856 n175__vdd n242__vdd 15.7583
rk2857 n177__vdd n243__vdd 15.7797
rk2858 n178__vdd n244__vdd 15.8451
rk2859 n178__vdd n245__vdd 15.8451
rk2860 n179__vdd n246__vdd 15.8665
rk2861 n179__vdd n247__vdd 15.8665
rk2862 n180__vdd n248__vdd 15.7761
rk2863 n180__vdd n249__vdd 15.7761
rk2864 n181__vdd n250__vdd 15.8539
rk2865 n181__vdd n251__vdd 15.8522
rk2866 n182__vdd n252__vdd 15.7671
rk2867 n183__vdd n253__vdd 15.7735
rk2868 n184__vdd n254__vdd 15.7797
rk2869 n185__vdd n255__vdd 15.7668
rk2870 n186__vdd n256__vdd 15.7882
rk2871 n187__vdd n257__vdd 15.7583
rk2872 n188__vdd n258__vdd 15.7627
rk2873 n189__vdd n259__vdd 15.7797
rk2874 n190__vdd n261__vdd 393e-3
rk2875 n261__vdd n262__vdd 75.4999
rk2876 n191__vdd n263__vdd 15.8814
rk2877 n191__vdd n264__vdd 15.8665
rk2878 n192__vdd n265__vdd 15.7583
rk2879 n193__vdd n266__vdd 15.7767
rk2880 n194__vdd n267__vdd 15.763
rk2881 n195__vdd n269__vdd 355.4e-3
rk2882 n269__vdd n270__vdd 75.4999
rk2883 n196__vdd n271__vdd 15.7583
rk2884 n198__vdd n272__vdd 15.8451
rk2885 n198__vdd n273__vdd 15.8451
rk2886 n199__vdd n274__vdd 15.8451
rk2887 n199__vdd n275__vdd 15.8451
rk2888 n200__vdd n276__vdd 15.8451
rk2889 n200__vdd n277__vdd 15.8451
rk2890 n201__vdd n278__vdd 15.8451
rk2891 n201__vdd n279__vdd 15.8451
rk2892 n202__vdd n280__vdd 62.4486
rk2893 n202__vdd n281__vdd 62.4486
rk2894 n203__vdd n282__vdd 62.4771
rk2895 n203__vdd n283__vdd 62.4771
rk2896 n205__vdd n284__vdd 15.8451
rk2897 n205__vdd n285__vdd 15.8451
rk2898 n206__vdd n286__vdd 15.8451
rk2899 n206__vdd n287__vdd 15.8451
rk2900 n207__vdd n288__vdd 62.5087
rk2901 n207__vdd n289__vdd 62.5087
rk2902 n209__vdd n290__vdd 31.2395
rk2903 n134__vdd n135__vdd 25
rk2904 n134__vdd n137__vdd 25
rk2905 n134__vdd n140__vdd 12.5
rk2906 n134__vdd n145__vdd 3.75
rk2907 n134__vdd n149__vdd 3.75
rk2908 n134__vdd n155__vdd 25
rk2909 n134__vdd n159__vdd 7.5
rk2910 n134__vdd n167__vdd 3.75
rk2911 n134__vdd n172__vdd 25
rk2912 n134__vdd n176__vdd 18.75
rk2913 n134__vdd n180__vdd 5.3571
rk2914 n134__vdd n188__vdd 3.75
rk2915 n134__vdd n197__vdd 3.75
rk2916 n134__vdd n204__vdd 3.75
rk2917 n134__vdd n208__vdd 3.75
rk2918 n260__vdd n261__vdd 31
rk2919 n268__vdd n269__vdd 31
rk2920 n291__vdd n292__vdd 31.4047
rk2921 n292__vdd n294__vdd 57.54e-3
rk2922 n294__vdd n295__vdd 33.07e-3
rk2923 n295__vdd n296__vdd 107.2e-3
rk2924 n296__vdd n297__vdd 23.5e-3
rk2925 n297__vdd n298__vdd 399.7e-3
rk2926 n298__vdd n299__vdd 25.66e-3
rk2927 n299__vdd n300__vdd 70.37e-3
rk2928 n300__vdd n301__vdd 53.41e-3
rk2929 n301__vdd n302__vdd 84.6e-3
rk2930 n302__vdd n303__vdd 96.04e-3
rk2931 n303__vdd n304__vdd 17.35e-3
rk2932 n304__vdd n305__vdd 36.06e-3
rk2933 n305__vdd n306__vdd 220.8e-3
rk2934 n306__vdd n307__vdd 84.6e-3
rk2935 n307__vdd n308__vdd 155.6e-3
rk2936 n308__vdd n309__vdd 75.57e-3
rk2937 n309__vdd n310__vdd 432.4e-3
rk2938 n310__vdd n311__vdd 855.6e-3
rk2939 n311__vdd n312__vdd 293e-3
rk2940 n312__vdd n313__vdd 64.39e-3
rk2941 n313__vdd n314__vdd 33.28e-3
rk2942 n314__vdd n315__vdd 109.8e-3
rk2943 n315__vdd n316__vdd 23.71e-3
rk2944 n316__vdd n317__vdd 124e-3
rk2945 n317__vdd n318__vdd 23.71e-3
rk2946 n318__vdd n319__vdd 109.8e-3
rk2947 n319__vdd n320__vdd 33.28e-3
rk2948 n320__vdd n321__vdd 64.39e-3
rk2949 n321__vdd n322__vdd 131.2e-3
rk2950 n322__vdd n323__vdd 33.28e-3
rk2951 n323__vdd n324__vdd 64.39e-3
rk2952 n324__vdd n325__vdd 804.5e-3
rk2953 n325__vdd n326__vdd 110.4e-3
rk2954 n326__vdd n327__vdd 35.46e-3
rk2955 n327__vdd n328__vdd 25.89e-3
rk2956 n328__vdd n329__vdd 97.25e-3
rk2957 n329__vdd n330__vdd 110.4e-3
rk2958 n330__vdd n331__vdd 61.36e-3
rk2959 n331__vdd n332__vdd 189.8e-3
rk2960 n332__vdd n333__vdd 64.18e-3
rk2961 n333__vdd n334__vdd 97.25e-3
rk2962 n334__vdd n335__vdd 265.9e-3
rk2963 n335__vdd n336__vdd 144.3e-3
rk2964 n336__vdd n337__vdd 168.3e-3
rk2965 n337__vdd n338__vdd 110.4e-3
rk2966 n338__vdd n339__vdd 61.36e-3
rk2967 n339__vdd n340__vdd 97.25e-3
rk2968 n340__vdd n341__vdd 110.4e-3
rk2969 n341__vdd n342__vdd 22.3e-3
rk2970 n342__vdd n343__vdd 39.05e-3
rk2971 n343__vdd n4__vdd 42.64e-3
rk2972 n4__vdd n344__vdd 211.3e-3
rk2973 n344__vdd n345__vdd 97.25e-3
rk2974 n345__vdd n346__vdd 181.4e-3
rk2975 n346__vdd n347__vdd 88.33e-3
rk2976 n347__vdd n348__vdd 62.4083
rk2977 n292__vdd n349__vdd 31.3477
rk2978 n295__vdd n350__vdd 31.4136
rk2979 n295__vdd n351__vdd 31.4136
rk2980 n297__vdd n352__vdd 31.4136
rk2981 n297__vdd n353__vdd 31.4136
rk2982 n298__vdd n354__vdd 15.8524
rk2983 n298__vdd n355__vdd 15.8524
rk2984 n300__vdd n356__vdd 15.8524
rk2985 n300__vdd n357__vdd 15.8524
rk2986 n301__vdd n358__vdd 15.8524
rk2987 n301__vdd n359__vdd 15.8524
rk2988 n302__vdd n360__vdd 15.8524
rk2989 n302__vdd n361__vdd 15.8524
rk2990 n303__vdd n362__vdd 62.4559
rk2991 n303__vdd n363__vdd 62.4559
rk2992 n305__vdd n364__vdd 62.4844
rk2993 n305__vdd n365__vdd 62.4844
rk2994 n306__vdd n366__vdd 15.8524
rk2995 n306__vdd n367__vdd 15.8524
rk2996 n307__vdd n368__vdd 15.8524
rk2997 n307__vdd n369__vdd 15.8524
rk2998 n309__vdd n370__vdd 62.5189
rk2999 n309__vdd n371__vdd 62.5189
rk3000 n310__vdd n372__vdd 15.7623
rk3001 n310__vdd n373__vdd 15.7623
rk3002 n311__vdd n374__vdd 31.2948
rk3003 n311__vdd n375__vdd 31.2948
rk3004 n312__vdd n376__vdd 15.7797
rk3005 n314__vdd n377__vdd 15.7583
rk3006 n316__vdd n378__vdd 31.3268
rk3007 n317__vdd n379__vdd 31.3268
rk3008 n319__vdd n380__vdd 31.3268
rk3009 n321__vdd n381__vdd 31.3375
rk3010 n322__vdd n382__vdd 15.7583
rk3011 n324__vdd n383__vdd 15.7797
rk3012 n325__vdd n384__vdd 15.8451
rk3013 n325__vdd n385__vdd 15.8451
rk3014 n326__vdd n386__vdd 15.8451
rk3015 n326__vdd n387__vdd 15.8451
rk3016 n328__vdd n388__vdd 15.8451
rk3017 n328__vdd n389__vdd 15.8451
rk3018 n329__vdd n390__vdd 15.8451
rk3019 n329__vdd n391__vdd 15.8451
rk3020 n330__vdd n392__vdd 62.4486
rk3021 n330__vdd n393__vdd 62.4486
rk3022 n331__vdd n394__vdd 62.4771
rk3023 n331__vdd n395__vdd 62.4771
rk3024 n333__vdd n396__vdd 15.8451
rk3025 n333__vdd n397__vdd 15.8451
rk3026 n334__vdd n398__vdd 15.8451
rk3027 n334__vdd n399__vdd 15.8451
rk3028 n335__vdd n400__vdd 62.5087
rk3029 n335__vdd n401__vdd 62.5087
rk3030 n337__vdd n402__vdd 15.8451
rk3031 n337__vdd n403__vdd 15.8451
rk3032 n338__vdd n404__vdd 15.8451
rk3033 n338__vdd n405__vdd 15.8451
rk3034 n339__vdd n406__vdd 15.8451
rk3035 n339__vdd n407__vdd 15.8451
rk3036 n340__vdd n408__vdd 15.8451
rk3037 n340__vdd n409__vdd 15.8451
rk3038 n341__vdd n410__vdd 62.4486
rk3039 n341__vdd n411__vdd 62.4486
rk3040 n343__vdd n412__vdd 62.4771
rk3041 n343__vdd n413__vdd 62.4771
rk3042 n344__vdd n414__vdd 15.8451
rk3043 n344__vdd n415__vdd 15.8451
rk3044 n345__vdd n416__vdd 15.8451
rk3045 n345__vdd n417__vdd 15.8451
rk3046 n347__vdd n418__vdd 62.5084
rk3047 n293__vdd n294__vdd 25
rk3048 n293__vdd n296__vdd 25
rk3049 n293__vdd n299__vdd 12.5
rk3050 n293__vdd n304__vdd 3.75
rk3051 n293__vdd n308__vdd 3.75
rk3052 n293__vdd n313__vdd 25
rk3053 n293__vdd n315__vdd 25
rk3054 n293__vdd n318__vdd 25
rk3055 n293__vdd n320__vdd 25
rk3056 n293__vdd n323__vdd 25
rk3057 n293__vdd n327__vdd 5.3571
rk3058 n293__vdd n332__vdd 3.75
rk3059 n293__vdd n336__vdd 3.75
rk3060 n293__vdd n342__vdd 3.75
rk3061 n293__vdd n346__vdd 3.75
rk3062 n4__serial_out_b_high_buff n5__serial_out_b_high_buff 640.9e-3
rk3063 n5__serial_out_b_high_buff n6__serial_out_b_high_buff 37.5134
rk3064 n5__serial_out_b_high_buff n7__serial_out_b_high_buff 13.1042
rk3065 n715__vss n716__vss 75.2804
rk3066 n716__vss n717__vss 57.54e-3
rk3067 n717__vss n718__vss 33.07e-3
rk3068 n718__vss n719__vss 107.2e-3
rk3069 n719__vss n720__vss 23.5e-3
rk3070 n720__vss n721__vss 399.7e-3
rk3071 n721__vss n722__vss 25.66e-3
rk3072 n722__vss n723__vss 70.37e-3
rk3073 n723__vss n724__vss 53.41e-3
rk3074 n724__vss n725__vss 84.6e-3
rk3075 n725__vss n726__vss 69e-3
rk3076 n726__vss n727__vss 44.38e-3
rk3077 n727__vss n728__vss 257.5e-3
rk3078 n728__vss n729__vss 84.6e-3
rk3079 n729__vss n730__vss 53.41e-3
rk3080 n730__vss n731__vss 101.6e-3
rk3081 n716__vss n732__vss 75.2196
rk3082 n718__vss n733__vss 75.2937
rk3083 n718__vss n734__vss 75.2937
rk3084 n720__vss n735__vss 75.2937
rk3085 n720__vss n736__vss 75.2937
rk3086 n721__vss n737__vss 37.7668
rk3087 n721__vss n738__vss 37.7668
rk3088 n723__vss n739__vss 37.7668
rk3089 n723__vss n740__vss 37.7668
rk3090 n724__vss n741__vss 37.7668
rk3091 n724__vss n742__vss 37.7668
rk3092 n725__vss n743__vss 37.7668
rk3093 n725__vss n744__vss 37.7668
rk3094 n726__vss n745__vss 75.2968
rk3095 n726__vss n746__vss 75.2968
rk3096 n728__vss n747__vss 37.7668
rk3097 n728__vss n748__vss 37.7668
rk3098 n729__vss n749__vss 37.7668
rk3099 n729__vss n750__vss 37.7668
rk3100 n730__vss n751__vss 75.3011
rk3101 n730__vss n752__vss 75.3011
rk3102 n731__vss n753__vss 75.1882
rk3103 n731__vss n754__vss 467.5e-3
rk3104 n754__vss n755__vss 37.7668
rk3105 n731__vss n756__vss 75.1882
rk3106 n754__vss n757__vss 374.3e-3
rk3107 n757__vss n758__vss 75.298
rk3108 n754__vss n759__vss 37.7668
rk3109 n757__vss n760__vss 148.9e-3
rk3110 n760__vss n761__vss 141.9e-3
rk3111 n761__vss n762__vss 37.6834
rk3112 n757__vss n763__vss 75.298
rk3113 n760__vss n764__vss 25.2316
rk3114 n761__vss n765__vss 17.73e-3
rk3115 n765__vss n766__vss 79.94e-3
rk3116 n766__vss n767__vss 37.6727
rk3117 n766__vss n768__vss 55.8e-3
rk3118 n768__vss n769__vss 53.62e-3
rk3119 n769__vss n770__vss 23.71e-3
rk3120 n770__vss n771__vss 75.207
rk3121 n768__vss n772__vss 37.6727
rk3122 n770__vss n773__vss 33.07e-3
rk3123 n773__vss n774__vss 61.78e-3
rk3124 n774__vss n775__vss 28.28e-3
rk3125 n775__vss n776__vss 75.207
rk3126 n773__vss n777__vss 37.6727
rk3127 n774__vss n778__vss 37.6727
rk3128 n775__vss n779__vss 23.71e-3
rk3129 n779__vss n780__vss 45.25e-3
rk3130 n780__vss n781__vss 64.17e-3
rk3131 n781__vss n782__vss 75.207
rk3132 n780__vss n783__vss 37.6727
rk3133 n781__vss n784__vss 15.12e-3
rk3134 n784__vss n785__vss 17.73e-3
rk3135 n785__vss n786__vss 64.39e-3
rk3136 n786__vss n787__vss 75.2123
rk3137 n784__vss n788__vss 75.2027
rk3138 n786__vss n789__vss 131.2e-3
rk3139 n789__vss n790__vss 37.6727
rk3140 n789__vss n791__vss 33.28e-3
rk3141 n791__vss n792__vss 64.39e-3
rk3142 n792__vss n793__vss 37.6834
rk3143 n792__vss n794__vss 35.46e-3
rk3144 n794__vss n795__vss 97.67e-3
rk3145 n795__vss n796__vss 61.78e-3
rk3146 n796__vss n797__vss 110.8e-3
rk3147 n797__vss n798__vss 252.2e-3
rk3148 n798__vss n799__vss 196e-3
rk3149 n799__vss n800__vss 48.62e-3
rk3150 n800__vss n801__vss 37.6727
rk3151 n794__vss n802__vss 37.6727
rk3152 n795__vss n803__vss 37.6727
rk3153 n796__vss n804__vss 75.207
rk3154 n797__vss n805__vss 75.2047
rk3155 n799__vss n806__vss 37.6727
rk3156 n800__vss n807__vss 48.62e-3
rk3157 n807__vss n808__vss 61.78e-3
rk3158 n808__vss n809__vss 37.6727
rk3159 n807__vss n810__vss 37.6834
rk3160 n808__vss n811__vss 35.68e-3
rk3161 n811__vss n812__vss 26.1e-3
rk3162 n812__vss n813__vss 37.6727
rk3163 n811__vss n814__vss 37.6798
rk3164 n812__vss n815__vss 71.35e-3
rk3165 n815__vss n816__vss 25.89e-3
rk3166 n816__vss n817__vss 37.6727
rk3167 n815__vss n818__vss 37.678
rk3168 n816__vss n819__vss 30.68e-3
rk3169 n819__vss n820__vss 48.62e-3
rk3170 n820__vss n821__vss 75.2027
rk3171 n819__vss n822__vss 37.678
rk3172 n820__vss n823__vss 48.62e-3
rk3173 n823__vss n824__vss 97.67e-3
rk3174 n824__vss n825__vss 97.67e-3
rk3175 n825__vss n826__vss 38.07e-3
rk3176 n826__vss n827__vss 24.91e-3
rk3177 n827__vss n828__vss 39.05e-3
rk3178 n828__vss n829__vss 37.6727
rk3179 n823__vss n830__vss 37.6834
rk3180 n824__vss n831__vss 37.6834
rk3181 n825__vss n832__vss 37.6727
rk3182 n827__vss n834__vss 205.2e-3
rk3183 n828__vss n403__vss 75.15e-3
rk3184 n403__vss n835__vss 22.52e-3
rk3185 n835__vss n836__vss 37.6727
rk3186 n834__vss n837__vss 31.3882
rk3187 n835__vss n838__vss 23.5e-3
rk3188 n838__vss n839__vss 37.85e-3
rk3189 n839__vss n840__vss 75.207
rk3190 n838__vss n841__vss 37.6848
rk3191 n839__vss n842__vss 109.1e-3
rk3192 n842__vss n843__vss 75.2099
rk3193 n842__vss n844__vss 12.22e-3
rk3194 n844__vss n845__vss 159.9e-3
rk3195 n845__vss n846__vss 66.78e-3
rk3196 n846__vss n847__vss 53.62e-3
rk3197 n847__vss n848__vss 112.2e-3
rk3198 n848__vss n849__vss 37.7411
rk3199 n844__vss n850__vss 37.6848
rk3200 n845__vss n852__vss 207e-3
rk3201 n852__vss n853__vss 31.3888
rk3202 n847__vss n854__vss 37.6727
rk3203 n848__vss n855__vss 59.57e-3
rk3204 n855__vss n856__vss 52.21e-3
rk3205 n856__vss n857__vss 37.6727
rk3206 n848__vss n858__vss 37.7437
rk3207 n855__vss n859__vss 37.6727
rk3208 n856__vss n860__vss 45.03e-3
rk3209 n860__vss n861__vss 16.32e-3
rk3210 n861__vss n862__vss 37.6727
rk3211 n860__vss n863__vss 37.6727
rk3212 n861__vss n864__vss 62.98e-3
rk3213 n864__vss n865__vss 34.27e-3
rk3214 n865__vss n866__vss 37.6727
rk3215 n864__vss n867__vss 75.2027
rk3216 n865__vss n868__vss 79.72e-3
rk3217 n868__vss n869__vss 75.2027
rk3218 n868__vss n870__vss 53.62e-3
rk3219 n870__vss n871__vss 179.2e-3
rk3220 n871__vss n872__vss 97.67e-3
rk3221 n872__vss n873__vss 16.32e-3
rk3222 n873__vss n874__vss 37.6727
rk3223 n871__vss n875__vss 37.6727
rk3224 n872__vss n876__vss 37.6727
rk3225 n873__vss n877__vss 45.03e-3
rk3226 n877__vss n878__vss 52.21e-3
rk3227 n878__vss n879__vss 37.6727
rk3228 n877__vss n880__vss 75.207
rk3229 n878__vss n881__vss 59.57e-3
rk3230 n881__vss n882__vss 75.2754
rk3231 n881__vss n883__vss 120.8e-3
rk3232 n883__vss n884__vss 75.2011
rk3233 n881__vss n885__vss 75.2757
rk3234 n883__vss n886__vss 75.3975
rk3235 n640__vss n717__vss 20.6667
rk3236 n640__vss n719__vss 20.6667
rk3237 n640__vss n722__vss 10.3333
rk3238 n640__vss n727__vss 3.1
rk3239 n640__vss n731__vss 3.1
rk3240 n640__vss n765__vss 10.3333
rk3241 n640__vss n769__vss 20.6667
rk3242 n640__vss n779__vss 20.6667
rk3243 n640__vss n785__vss 20.6667
rk3244 n640__vss n791__vss 20.6667
rk3245 n640__vss n798__vss 20.6667
rk3246 n640__vss n811__vss 4.4286
rk3247 n640__vss n826__vss 3.1
rk3248 n833__vss n834__vss 75
rk3249 n640__vss n846__vss 3.1
rk3250 n851__vss n852__vss 75
rk3251 n640__vss n870__vss 3.1
rk3252 n640__vss n883__vss 3.1
rk3253 n887__vss n888__vss 75.2838
rk3254 n888__vss n889__vss 33.28e-3
rk3255 n889__vss n890__vss 107.5e-3
rk3256 n890__vss n891__vss 23.71e-3
rk3257 n891__vss n892__vss 404.7e-3
rk3258 n892__vss n893__vss 81.02e-3
rk3259 n893__vss n894__vss 22.06e-3
rk3260 n894__vss n895__vss 57.47e-3
rk3261 n895__vss n896__vss 90.84e-3
rk3262 n896__vss n897__vss 74.16e-3
rk3263 n897__vss n898__vss 154.4e-3
rk3264 n898__vss n899__vss 168.9e-3
rk3265 n899__vss n900__vss 35.22e-3
rk3266 n900__vss n901__vss 55.25e-3
rk3267 n901__vss n902__vss 59.71e-3
rk3268 n902__vss n903__vss 100.9e-3
rk3269 n903__vss n904__vss 49.68e-3
rk3270 n904__vss n905__vss 62.11e-3
rk3271 n905__vss n906__vss 393.6e-3
rk3272 n906__vss n907__vss 24.1e-3
rk3273 n907__vss n908__vss 120.6e-3
rk3274 n908__vss n530__vss 138.8e-3
rk3275 n530__vss n909__vss 23.71e-3
rk3276 n909__vss n910__vss 71.35e-3
rk3277 n910__vss n911__vss 339.5e-3
rk3278 n911__vss n912__vss 105.1e-3
rk3279 n912__vss n913__vss 126.4e-3
rk3280 n913__vss n914__vss 159.9e-3
rk3281 n914__vss n503__vss 88.67e-3
rk3282 n503__vss n915__vss 79.31e-3
rk3283 n915__vss n916__vss 334.7e-3
rk3284 n916__vss n917__vss 239e-3
rk3285 n917__vss n918__vss 277.3e-3
rk3286 n918__vss n919__vss 148.9e-3
rk3287 n919__vss n920__vss 110.4e-3
rk3288 n920__vss n921__vss 35.46e-3
rk3289 n921__vss n922__vss 25.89e-3
rk3290 n922__vss n923__vss 97.25e-3
rk3291 n923__vss n924__vss 79.3e-3
rk3292 n924__vss n925__vss 283.1e-3
rk3293 n925__vss n926__vss 64.18e-3
rk3294 n926__vss n406__vss 74.94e-3
rk3295 n406__vss n927__vss 22.3e-3
rk3296 n927__vss n928__vss 61.36e-3
rk3297 n928__vss n929__vss 110.4e-3
rk3298 n929__vss n930__vss 237.6e-3
rk3299 n930__vss n931__vss 168.3e-3
rk3300 n931__vss n932__vss 110.4e-3
rk3301 n932__vss n933__vss 61.36e-3
rk3302 n933__vss n934__vss 97.25e-3
rk3303 n934__vss n935__vss 79.3e-3
rk3304 n935__vss n936__vss 53.41e-3
rk3305 n936__vss n937__vss 293.9e-3
rk3306 n937__vss n938__vss 97.25e-3
rk3307 n938__vss n939__vss 61.36e-3
rk3308 n939__vss n940__vss 119.2e-3
rk3309 n889__vss n941__vss 75.207
rk3310 n891__vss n942__vss 75.207
rk3311 n892__vss n943__vss 37.6743
rk3312 n894__vss n944__vss 37.6743
rk3313 n895__vss n945__vss 37.6743
rk3314 n896__vss n946__vss 37.6743
rk3315 n897__vss n947__vss 75.2042
rk3316 n899__vss n948__vss 37.6743
rk3317 n900__vss n949__vss 75.1957
rk3318 n901__vss n950__vss 37.6743
rk3319 n902__vss n951__vss 75.3218
rk3320 n902__vss n952__vss 75.3297
rk3321 n903__vss n953__vss 75.2063
rk3322 n904__vss n954__vss 37.6614
rk3323 n906__vss n955__vss 37.6743
rk3324 n907__vss n956__vss 75.1957
rk3325 n908__vss n957__vss 75.2216
rk3326 n909__vss n958__vss 37.6727
rk3327 n910__vss n959__vss 75.2112
rk3328 n912__vss n960__vss 75.207
rk3329 n913__vss n961__vss 75.212
rk3330 n914__vss n962__vss 37.6727
rk3331 n916__vss n963__vss 75.207
rk3332 n918__vss n964__vss 75.207
rk3333 n919__vss n965__vss 37.7595
rk3334 n919__vss n966__vss 37.7595
rk3335 n920__vss n967__vss 37.7595
rk3336 n920__vss n968__vss 37.7595
rk3337 n922__vss n969__vss 37.7595
rk3338 n922__vss n970__vss 37.7595
rk3339 n923__vss n971__vss 37.7595
rk3340 n923__vss n972__vss 37.7595
rk3341 n924__vss n973__vss 75.2895
rk3342 n924__vss n974__vss 75.2895
rk3343 n926__vss n975__vss 37.7595
rk3344 n926__vss n976__vss 37.7595
rk3345 n927__vss n977__vss 37.7595
rk3346 n927__vss n978__vss 37.7595
rk3347 n928__vss n979__vss 75.2937
rk3348 n928__vss n980__vss 75.2937
rk3349 n929__vss n981__vss 75.2915
rk3350 n929__vss n982__vss 75.2915
rk3351 n931__vss n983__vss 37.7595
rk3352 n931__vss n984__vss 37.7595
rk3353 n932__vss n985__vss 37.7595
rk3354 n932__vss n986__vss 37.7595
rk3355 n933__vss n987__vss 37.7595
rk3356 n933__vss n988__vss 37.7595
rk3357 n934__vss n989__vss 37.7595
rk3358 n934__vss n990__vss 37.7595
rk3359 n935__vss n991__vss 75.2895
rk3360 n935__vss n992__vss 75.2895
rk3361 n937__vss n993__vss 37.7595
rk3362 n937__vss n994__vss 37.7595
rk3363 n938__vss n995__vss 37.7595
rk3364 n938__vss n996__vss 37.7595
rk3365 n939__vss n997__vss 75.2937
rk3366 n939__vss n998__vss 75.2937
rk3367 n940__vss n999__vss 75.2011
rk3368 n940__vss n1000__vss 75.2011
rk3369 n640__vss n888__vss 20.6667
rk3370 n640__vss n890__vss 20.6667
rk3371 n640__vss n893__vss 6.2
rk3372 n640__vss n898__vss 3.1
rk3373 n640__vss n905__vss 3.1
rk3374 n640__vss n908__vss 3.1
rk3375 n640__vss n911__vss 3.1
rk3376 n640__vss n915__vss 3.1
rk3377 n640__vss n917__vss 3.1
rk3378 n640__vss n921__vss 4.4286
rk3379 n640__vss n925__vss 3.1
rk3380 n640__vss n930__vss 3.1
rk3381 n640__vss n936__vss 3.1
rk3382 n640__vss n940__vss 3.1
rk3383 n1001__vss n1002__vss 10.7834
rk3384 n1002__vss n1003__vss 644.2e-3
rk3385 n1003__vss n1004__vss 6.1924
rk3386 n1002__vss n1005__vss 5.5602
rk3387 n678__vddio n679__vddio 7.1062
rk3388 n679__vddio n680__vddio 847e-3
rk3389 n680__vddio n681__vddio 4.4452
rk3390 n679__vddio n682__vddio 3.6209
rk3391 n8__serial_out_b_high_buff n2__serial_out_b_high_buff 23.0122
rk3392 n683__vddio n684__vddio 25.2185
rk3393 n684__vddio n685__vddio 12.8226
rk3394 n687__vddio n688__vddio 84.92e-3
rk3395 n688__vddio n689__vddio 327.8e-3
rk3396 n689__vddio n690__vddio 574.2e-3
rk3397 n690__vddio n691__vddio 574.2e-3
rk3398 n691__vddio n692__vddio 574.2e-3
rk3399 n692__vddio n693__vddio 574.2e-3
rk3400 n693__vddio n694__vddio 574.2e-3
rk3401 n694__vddio n695__vddio 574.2e-3
rk3402 n695__vddio n696__vddio 574.2e-3
rk3403 n696__vddio n417__vddio 447.4e-3
rk3404 n417__vddio n697__vddio 126.8e-3
rk3405 n697__vddio n698__vddio 41.66e-3
rk3406 n698__vddio n407__vddio 441.3e-3
rk3407 n407__vddio n700__vddio 527.6e-3
rk3408 n698__vddio n701__vddio 164.7e-3
rk3409 n701__vddio n702__vddio 167.1e-3
rk3410 n702__vddio n703__vddio 167.1e-3
rk3411 n703__vddio n704__vddio 32.09e-3
rk3412 n704__vddio n705__vddio 135e-3
rk3413 n705__vddio n706__vddio 167.1e-3
rk3414 n706__vddio n707__vddio 167.1e-3
rk3415 n707__vddio n708__vddio 103.9e-3
rk3416 n708__vddio n709__vddio 63.19e-3
rk3417 n709__vddio n710__vddio 167.1e-3
rk3418 n710__vddio n711__vddio 167.1e-3
rk3419 n711__vddio n712__vddio 175.6e-3
rk3420 n712__vddio n713__vddio 158.9e-3
rk3421 n713__vddio n714__vddio 167.1e-3
rk3422 n714__vddio n715__vddio 167.1e-3
rk3423 n715__vddio n716__vddio 79.94e-3
rk3424 n716__vddio n717__vddio 87.12e-3
rk3425 n717__vddio n718__vddio 167.1e-3
rk3426 n718__vddio n719__vddio 167.1e-3
rk3427 n719__vddio n720__vddio 151.7e-3
rk3428 n720__vddio n721__vddio 15.34e-3
rk3429 n721__vddio n722__vddio 167.1e-3
rk3430 n722__vddio n723__vddio 167.1e-3
rk3431 n723__vddio n724__vddio 167.1e-3
rk3432 n724__vddio n725__vddio 56.01e-3
rk3433 n725__vddio n726__vddio 111e-3
rk3434 n726__vddio n727__vddio 167.1e-3
rk3435 n727__vddio n728__vddio 167.1e-3
rk3436 n728__vddio n729__vddio 127.8e-3
rk3437 n729__vddio n730__vddio 39.26e-3
rk3438 n730__vddio n731__vddio 167.1e-3
rk3439 n731__vddio n732__vddio 167.1e-3
rk3440 n732__vddio n733__vddio 167.1e-3
rk3441 n733__vddio n734__vddio 32.09e-3
rk3442 n734__vddio n735__vddio 135e-3
rk3443 n735__vddio n736__vddio 167.1e-3
rk3444 n736__vddio n737__vddio 167.1e-3
rk3445 n737__vddio n738__vddio 103.9e-3
rk3446 n738__vddio n739__vddio 63.19e-3
rk3447 n739__vddio n740__vddio 167.1e-3
rk3448 n740__vddio n741__vddio 167.1e-3
rk3449 n741__vddio n742__vddio 175.6e-3
rk3450 n742__vddio n743__vddio 158.9e-3
rk3451 n743__vddio n744__vddio 167.1e-3
rk3452 n744__vddio n745__vddio 167.1e-3
rk3453 n745__vddio n746__vddio 79.94e-3
rk3454 n746__vddio n747__vddio 87.12e-3
rk3455 n747__vddio n748__vddio 167.1e-3
rk3456 n748__vddio n749__vddio 167.1e-3
rk3457 n749__vddio n750__vddio 151.7e-3
rk3458 n750__vddio n751__vddio 15.34e-3
rk3459 n751__vddio n752__vddio 167.1e-3
rk3460 n752__vddio n753__vddio 167.1e-3
rk3461 n753__vddio n754__vddio 167.1e-3
rk3462 n754__vddio n755__vddio 56.01e-3
rk3463 n755__vddio n756__vddio 111e-3
rk3464 n756__vddio n757__vddio 167.1e-3
rk3465 n757__vddio n758__vddio 167.1e-3
rk3466 n758__vddio n759__vddio 127.8e-3
rk3467 n759__vddio n760__vddio 39.26e-3
rk3468 n760__vddio n761__vddio 167.1e-3
rk3469 n761__vddio n7__vddio 599.6e-3
rk3470 n7__vddio n763__vddio 528.5e-3
rk3471 n763__vddio n6__vddio 116e-3
rk3472 n6__vddio n3__vddio 1.1789
rk3473 n3__vddio n764__vddio 201e-3
rk3474 n764__vddio n2__vddio 1.0839
rk3475 n2__vddio n765__vddio 441.8e-3
rk3476 n765__vddio n762__vddio 8.8496
rk3477 n700__vddio n406__vddio 111.9e-3
rk3478 n406__vddio n403__vddio 1.1771
rk3479 n403__vddio n766__vddio 200.1e-3
rk3480 n766__vddio n402__vddio 1.083
rk3481 n402__vddio n767__vddio 440.9e-3
rk3482 n767__vddio n699__vddio 8.8496
rk3483 n701__vddio n399__vddio 438e-3
rk3484 n399__vddio n769__vddio 524.2e-3
rk3485 n769__vddio n398__vddio 104.4e-3
rk3486 n398__vddio n395__vddio 1.1705
rk3487 n395__vddio n770__vddio 196.8e-3
rk3488 n770__vddio n394__vddio 1.0796
rk3489 n394__vddio n771__vddio 437.6e-3
rk3490 n771__vddio n768__vddio 8.8496
rk3491 n702__vddio n392__vddio 438e-3
rk3492 n392__vddio n773__vddio 524.2e-3
rk3493 n773__vddio n389__vddio 104.4e-3
rk3494 n389__vddio n388__vddio 1.1705
rk3495 n388__vddio n774__vddio 196.8e-3
rk3496 n774__vddio n385__vddio 1.0796
rk3497 n385__vddio n775__vddio 437.6e-3
rk3498 n775__vddio n772__vddio 8.8496
rk3499 n703__vddio n383__vddio 441.3e-3
rk3500 n383__vddio n777__vddio 527.6e-3
rk3501 n777__vddio n382__vddio 111.9e-3
rk3502 n382__vddio n379__vddio 1.1771
rk3503 n379__vddio n778__vddio 200.1e-3
rk3504 n778__vddio n378__vddio 1.083
rk3505 n378__vddio n779__vddio 440.9e-3
rk3506 n779__vddio n776__vddio 8.8496
rk3507 n705__vddio n375__vddio 441.3e-3
rk3508 n375__vddio n781__vddio 527.6e-3
rk3509 n781__vddio n374__vddio 111.9e-3
rk3510 n374__vddio n371__vddio 1.1771
rk3511 n371__vddio n782__vddio 200.1e-3
rk3512 n782__vddio n370__vddio 1.083
rk3513 n370__vddio n783__vddio 440.9e-3
rk3514 n783__vddio n780__vddio 8.8496
rk3515 n706__vddio n367__vddio 441.3e-3
rk3516 n367__vddio n785__vddio 527.6e-3
rk3517 n785__vddio n366__vddio 111.9e-3
rk3518 n366__vddio n363__vddio 1.1771
rk3519 n363__vddio n786__vddio 200.1e-3
rk3520 n786__vddio n362__vddio 1.083
rk3521 n362__vddio n787__vddio 440.9e-3
rk3522 n787__vddio n784__vddio 8.8496
rk3523 n707__vddio n359__vddio 441.3e-3
rk3524 n359__vddio n789__vddio 527.6e-3
rk3525 n789__vddio n358__vddio 111.9e-3
rk3526 n358__vddio n355__vddio 1.1771
rk3527 n355__vddio n790__vddio 200.1e-3
rk3528 n790__vddio n354__vddio 1.083
rk3529 n354__vddio n791__vddio 440.9e-3
rk3530 n791__vddio n788__vddio 8.8496
rk3531 n709__vddio n352__vddio 444.1e-3
rk3532 n352__vddio n793__vddio 530.3e-3
rk3533 n793__vddio n349__vddio 116e-3
rk3534 n349__vddio n348__vddio 1.1827
rk3535 n348__vddio n794__vddio 202.9e-3
rk3536 n794__vddio n345__vddio 1.0857
rk3537 n345__vddio n795__vddio 443.7e-3
rk3538 n795__vddio n792__vddio 8.8496
rk3539 n710__vddio n343__vddio 444.1e-3
rk3540 n343__vddio n797__vddio 530.3e-3
rk3541 n797__vddio n342__vddio 116e-3
rk3542 n342__vddio n339__vddio 1.1827
rk3543 n339__vddio n798__vddio 202.9e-3
rk3544 n798__vddio n338__vddio 1.0857
rk3545 n338__vddio n799__vddio 443.7e-3
rk3546 n799__vddio n796__vddio 8.8496
rk3547 n711__vddio n335__vddio 437.1e-3
rk3548 n335__vddio n801__vddio 523.4e-3
rk3549 n801__vddio n334__vddio 102.1e-3
rk3550 n334__vddio n331__vddio 1.1688
rk3551 n331__vddio n802__vddio 195.9e-3
rk3552 n802__vddio n330__vddio 1.0788
rk3553 n330__vddio n803__vddio 436.7e-3
rk3554 n803__vddio n800__vddio 8.8496
rk3555 n712__vddio n327__vddio 433.5e-3
rk3556 n327__vddio n805__vddio 523.4e-3
rk3557 n805__vddio n326__vddio 102.1e-3
rk3558 n326__vddio n323__vddio 1.1688
rk3559 n323__vddio n806__vddio 195.9e-3
rk3560 n806__vddio n322__vddio 1.0788
rk3561 n322__vddio n807__vddio 436.7e-3
rk3562 n807__vddio n804__vddio 8.8496
rk3563 n713__vddio n319__vddio 444.1e-3
rk3564 n319__vddio n809__vddio 530.3e-3
rk3565 n809__vddio n318__vddio 116e-3
rk3566 n318__vddio n315__vddio 1.1827
rk3567 n315__vddio n810__vddio 202.9e-3
rk3568 n810__vddio n314__vddio 1.0857
rk3569 n314__vddio n811__vddio 443.7e-3
rk3570 n811__vddio n808__vddio 8.8496
rk3571 n714__vddio n311__vddio 444.1e-3
rk3572 n311__vddio n813__vddio 530.3e-3
rk3573 n813__vddio n310__vddio 116e-3
rk3574 n310__vddio n307__vddio 1.1827
rk3575 n307__vddio n814__vddio 202.9e-3
rk3576 n814__vddio n306__vddio 1.0857
rk3577 n306__vddio n815__vddio 443.7e-3
rk3578 n815__vddio n812__vddio 8.8496
rk3579 n715__vddio n303__vddio 441.3e-3
rk3580 n303__vddio n817__vddio 527.6e-3
rk3581 n817__vddio n302__vddio 111.9e-3
rk3582 n302__vddio n299__vddio 1.1771
rk3583 n299__vddio n818__vddio 200.1e-3
rk3584 n818__vddio n298__vddio 1.083
rk3585 n298__vddio n819__vddio 440.9e-3
rk3586 n819__vddio n816__vddio 8.8496
rk3587 n717__vddio n295__vddio 441.3e-3
rk3588 n295__vddio n821__vddio 527.6e-3
rk3589 n821__vddio n294__vddio 111.9e-3
rk3590 n294__vddio n291__vddio 1.1771
rk3591 n291__vddio n822__vddio 200.1e-3
rk3592 n822__vddio n290__vddio 1.083
rk3593 n290__vddio n823__vddio 440.9e-3
rk3594 n823__vddio n820__vddio 8.8496
rk3595 n718__vddio n287__vddio 444.1e-3
rk3596 n287__vddio n825__vddio 530.3e-3
rk3597 n825__vddio n286__vddio 116e-3
rk3598 n286__vddio n283__vddio 1.1827
rk3599 n283__vddio n826__vddio 202.9e-3
rk3600 n826__vddio n282__vddio 1.0857
rk3601 n282__vddio n827__vddio 443.7e-3
rk3602 n827__vddio n824__vddio 8.8496
rk3603 n719__vddio n279__vddio 444.1e-3
rk3604 n279__vddio n829__vddio 530.3e-3
rk3605 n829__vddio n278__vddio 116e-3
rk3606 n278__vddio n275__vddio 1.1827
rk3607 n275__vddio n830__vddio 202.9e-3
rk3608 n830__vddio n274__vddio 1.0857
rk3609 n274__vddio n831__vddio 443.7e-3
rk3610 n831__vddio n828__vddio 8.8496
rk3611 n721__vddio n271__vddio 437.1e-3
rk3612 n271__vddio n833__vddio 523.4e-3
rk3613 n833__vddio n270__vddio 102.1e-3
rk3614 n270__vddio n267__vddio 1.1688
rk3615 n267__vddio n834__vddio 195.9e-3
rk3616 n834__vddio n266__vddio 1.0788
rk3617 n266__vddio n835__vddio 436.7e-3
rk3618 n835__vddio n832__vddio 8.8496
rk3619 n722__vddio n263__vddio 437.1e-3
rk3620 n263__vddio n837__vddio 523.4e-3
rk3621 n837__vddio n262__vddio 102.1e-3
rk3622 n262__vddio n259__vddio 1.1688
rk3623 n259__vddio n838__vddio 195.9e-3
rk3624 n838__vddio n258__vddio 1.0788
rk3625 n258__vddio n839__vddio 436.7e-3
rk3626 n839__vddio n836__vddio 8.8496
rk3627 n723__vddio n255__vddio 444.1e-3
rk3628 n255__vddio n841__vddio 530.3e-3
rk3629 n841__vddio n254__vddio 116e-3
rk3630 n254__vddio n251__vddio 1.1827
rk3631 n251__vddio n842__vddio 202.9e-3
rk3632 n842__vddio n250__vddio 1.0857
rk3633 n250__vddio n843__vddio 443.7e-3
rk3634 n843__vddio n840__vddio 8.8496
rk3635 n724__vddio n247__vddio 441.3e-3
rk3636 n247__vddio n845__vddio 527.6e-3
rk3637 n845__vddio n246__vddio 111.9e-3
rk3638 n246__vddio n243__vddio 1.1771
rk3639 n243__vddio n846__vddio 200.1e-3
rk3640 n846__vddio n242__vddio 1.083
rk3641 n242__vddio n847__vddio 440.9e-3
rk3642 n847__vddio n844__vddio 8.8496
rk3643 n726__vddio n239__vddio 441.3e-3
rk3644 n239__vddio n849__vddio 527.6e-3
rk3645 n849__vddio n238__vddio 111.9e-3
rk3646 n238__vddio n235__vddio 1.1771
rk3647 n235__vddio n850__vddio 200.1e-3
rk3648 n850__vddio n234__vddio 1.083
rk3649 n234__vddio n851__vddio 440.9e-3
rk3650 n851__vddio n848__vddio 8.8496
rk3651 n727__vddio n231__vddio 444.1e-3
rk3652 n231__vddio n853__vddio 530.3e-3
rk3653 n853__vddio n230__vddio 116e-3
rk3654 n230__vddio n227__vddio 1.1827
rk3655 n227__vddio n854__vddio 202.9e-3
rk3656 n854__vddio n226__vddio 1.0857
rk3657 n226__vddio n855__vddio 443.7e-3
rk3658 n855__vddio n852__vddio 8.8496
rk3659 n728__vddio n223__vddio 444.1e-3
rk3660 n223__vddio n857__vddio 530.3e-3
rk3661 n857__vddio n222__vddio 116e-3
rk3662 n222__vddio n219__vddio 1.1827
rk3663 n219__vddio n858__vddio 202.9e-3
rk3664 n858__vddio n218__vddio 1.0857
rk3665 n218__vddio n859__vddio 443.7e-3
rk3666 n859__vddio n856__vddio 8.8496
rk3667 n730__vddio n215__vddio 437.1e-3
rk3668 n215__vddio n861__vddio 523.4e-3
rk3669 n861__vddio n214__vddio 102.1e-3
rk3670 n214__vddio n211__vddio 1.1688
rk3671 n211__vddio n862__vddio 195.9e-3
rk3672 n862__vddio n210__vddio 1.0788
rk3673 n210__vddio n863__vddio 436.7e-3
rk3674 n863__vddio n860__vddio 8.8496
rk3675 n731__vddio n207__vddio 437.1e-3
rk3676 n207__vddio n865__vddio 523.4e-3
rk3677 n865__vddio n206__vddio 102.1e-3
rk3678 n206__vddio n203__vddio 1.1688
rk3679 n203__vddio n866__vddio 195.9e-3
rk3680 n866__vddio n202__vddio 1.0788
rk3681 n202__vddio n867__vddio 436.7e-3
rk3682 n867__vddio n864__vddio 8.8496
rk3683 n732__vddio n199__vddio 444.1e-3
rk3684 n199__vddio n869__vddio 530.3e-3
rk3685 n869__vddio n198__vddio 116e-3
rk3686 n198__vddio n195__vddio 1.1827
rk3687 n195__vddio n870__vddio 202.9e-3
rk3688 n870__vddio n194__vddio 1.0857
rk3689 n194__vddio n871__vddio 443.7e-3
rk3690 n871__vddio n868__vddio 8.8496
rk3691 n733__vddio n191__vddio 444.1e-3
rk3692 n191__vddio n873__vddio 530.3e-3
rk3693 n873__vddio n190__vddio 116e-3
rk3694 n190__vddio n187__vddio 1.1827
rk3695 n187__vddio n874__vddio 202.9e-3
rk3696 n874__vddio n186__vddio 1.0857
rk3697 n186__vddio n875__vddio 443.7e-3
rk3698 n875__vddio n872__vddio 8.8496
rk3699 n735__vddio n183__vddio 441.3e-3
rk3700 n183__vddio n877__vddio 527.6e-3
rk3701 n877__vddio n182__vddio 111.9e-3
rk3702 n182__vddio n179__vddio 1.1771
rk3703 n179__vddio n878__vddio 200.1e-3
rk3704 n878__vddio n178__vddio 1.083
rk3705 n178__vddio n879__vddio 440.9e-3
rk3706 n879__vddio n876__vddio 8.8496
rk3707 n736__vddio n175__vddio 441.3e-3
rk3708 n175__vddio n881__vddio 527.6e-3
rk3709 n881__vddio n174__vddio 111.9e-3
rk3710 n174__vddio n171__vddio 1.1771
rk3711 n171__vddio n882__vddio 200.1e-3
rk3712 n882__vddio n170__vddio 1.083
rk3713 n170__vddio n883__vddio 440.9e-3
rk3714 n883__vddio n880__vddio 8.8496
rk3715 n737__vddio n167__vddio 444.1e-3
rk3716 n167__vddio n885__vddio 530.3e-3
rk3717 n885__vddio n166__vddio 116e-3
rk3718 n166__vddio n163__vddio 1.1827
rk3719 n163__vddio n886__vddio 202.9e-3
rk3720 n886__vddio n162__vddio 1.0857
rk3721 n162__vddio n887__vddio 443.7e-3
rk3722 n887__vddio n884__vddio 8.8496
rk3723 n739__vddio n159__vddio 444.1e-3
rk3724 n159__vddio n889__vddio 530.3e-3
rk3725 n889__vddio n158__vddio 116e-3
rk3726 n158__vddio n155__vddio 1.1827
rk3727 n155__vddio n890__vddio 202.9e-3
rk3728 n890__vddio n154__vddio 1.0857
rk3729 n154__vddio n891__vddio 443.7e-3
rk3730 n891__vddio n888__vddio 8.8496
rk3731 n740__vddio n151__vddio 437.1e-3
rk3732 n151__vddio n893__vddio 523.4e-3
rk3733 n893__vddio n150__vddio 102.1e-3
rk3734 n150__vddio n147__vddio 1.1688
rk3735 n147__vddio n894__vddio 195.9e-3
rk3736 n894__vddio n146__vddio 1.0788
rk3737 n146__vddio n895__vddio 436.7e-3
rk3738 n895__vddio n892__vddio 8.8496
rk3739 n741__vddio n143__vddio 437.1e-3
rk3740 n143__vddio n897__vddio 523.4e-3
rk3741 n897__vddio n142__vddio 102.1e-3
rk3742 n142__vddio n139__vddio 1.1688
rk3743 n139__vddio n898__vddio 195.9e-3
rk3744 n898__vddio n138__vddio 1.0788
rk3745 n138__vddio n899__vddio 436.7e-3
rk3746 n899__vddio n896__vddio 8.8496
rk3747 n742__vddio n135__vddio 440.4e-3
rk3748 n135__vddio n901__vddio 530.3e-3
rk3749 n901__vddio n134__vddio 116e-3
rk3750 n134__vddio n131__vddio 1.1827
rk3751 n131__vddio n902__vddio 202.9e-3
rk3752 n902__vddio n130__vddio 1.0857
rk3753 n130__vddio n903__vddio 443.7e-3
rk3754 n903__vddio n900__vddio 8.8496
rk3755 n743__vddio n127__vddio 442.2e-3
rk3756 n127__vddio n905__vddio 528.5e-3
rk3757 n905__vddio n126__vddio 116e-3
rk3758 n126__vddio n123__vddio 1.1789
rk3759 n123__vddio n906__vddio 201e-3
rk3760 n906__vddio n122__vddio 1.0839
rk3761 n122__vddio n907__vddio 441.8e-3
rk3762 n907__vddio n904__vddio 8.8496
rk3763 n744__vddio n119__vddio 442.2e-3
rk3764 n119__vddio n909__vddio 528.5e-3
rk3765 n909__vddio n118__vddio 116e-3
rk3766 n118__vddio n115__vddio 1.1789
rk3767 n115__vddio n910__vddio 201e-3
rk3768 n910__vddio n114__vddio 1.0839
rk3769 n114__vddio n911__vddio 441.8e-3
rk3770 n911__vddio n908__vddio 8.8496
rk3771 n745__vddio n111__vddio 438e-3
rk3772 n111__vddio n913__vddio 524.2e-3
rk3773 n913__vddio n110__vddio 104.4e-3
rk3774 n110__vddio n107__vddio 1.1705
rk3775 n107__vddio n914__vddio 196.8e-3
rk3776 n914__vddio n106__vddio 1.0796
rk3777 n106__vddio n915__vddio 437.6e-3
rk3778 n915__vddio n912__vddio 8.8496
rk3779 n747__vddio n103__vddio 438e-3
rk3780 n103__vddio n917__vddio 524.2e-3
rk3781 n917__vddio n102__vddio 104.4e-3
rk3782 n102__vddio n99__vddio 1.1705
rk3783 n99__vddio n918__vddio 196.8e-3
rk3784 n918__vddio n98__vddio 1.0796
rk3785 n98__vddio n919__vddio 437.6e-3
rk3786 n919__vddio n916__vddio 8.8496
rk3787 n748__vddio n95__vddio 441.3e-3
rk3788 n95__vddio n921__vddio 527.6e-3
rk3789 n921__vddio n94__vddio 111.9e-3
rk3790 n94__vddio n91__vddio 1.1771
rk3791 n91__vddio n922__vddio 200.1e-3
rk3792 n922__vddio n90__vddio 1.083
rk3793 n90__vddio n923__vddio 440.9e-3
rk3794 n923__vddio n920__vddio 8.8496
rk3795 n749__vddio n87__vddio 441.3e-3
rk3796 n87__vddio n925__vddio 527.6e-3
rk3797 n925__vddio n86__vddio 111.9e-3
rk3798 n86__vddio n83__vddio 1.1771
rk3799 n83__vddio n926__vddio 200.1e-3
rk3800 n926__vddio n82__vddio 1.083
rk3801 n82__vddio n927__vddio 440.9e-3
rk3802 n927__vddio n924__vddio 8.8496
rk3803 n751__vddio n79__vddio 444.1e-3
rk3804 n79__vddio n929__vddio 530.3e-3
rk3805 n929__vddio n78__vddio 116e-3
rk3806 n78__vddio n75__vddio 1.1827
rk3807 n75__vddio n930__vddio 202.9e-3
rk3808 n930__vddio n74__vddio 1.0857
rk3809 n74__vddio n931__vddio 443.7e-3
rk3810 n931__vddio n928__vddio 8.8496
rk3811 n752__vddio n71__vddio 444.1e-3
rk3812 n71__vddio n933__vddio 530.3e-3
rk3813 n933__vddio n70__vddio 116e-3
rk3814 n70__vddio n67__vddio 1.1827
rk3815 n67__vddio n934__vddio 202.9e-3
rk3816 n934__vddio n66__vddio 1.0857
rk3817 n66__vddio n935__vddio 443.7e-3
rk3818 n935__vddio n932__vddio 8.8496
rk3819 n753__vddio n63__vddio 442.2e-3
rk3820 n63__vddio n937__vddio 528.5e-3
rk3821 n937__vddio n62__vddio 116e-3
rk3822 n62__vddio n59__vddio 1.1789
rk3823 n59__vddio n938__vddio 201e-3
rk3824 n938__vddio n58__vddio 1.0839
rk3825 n58__vddio n939__vddio 441.8e-3
rk3826 n939__vddio n936__vddio 8.8496
rk3827 n754__vddio n55__vddio 442.2e-3
rk3828 n55__vddio n941__vddio 528.5e-3
rk3829 n941__vddio n54__vddio 116e-3
rk3830 n54__vddio n51__vddio 1.1789
rk3831 n51__vddio n942__vddio 201e-3
rk3832 n942__vddio n50__vddio 1.0839
rk3833 n50__vddio n943__vddio 441.8e-3
rk3834 n943__vddio n940__vddio 8.8496
rk3835 n756__vddio n47__vddio 438e-3
rk3836 n47__vddio n945__vddio 524.2e-3
rk3837 n945__vddio n46__vddio 104.4e-3
rk3838 n46__vddio n43__vddio 1.1705
rk3839 n43__vddio n946__vddio 196.8e-3
rk3840 n946__vddio n42__vddio 1.0796
rk3841 n42__vddio n947__vddio 437.6e-3
rk3842 n947__vddio n944__vddio 8.8496
rk3843 n757__vddio n39__vddio 438e-3
rk3844 n39__vddio n949__vddio 524.2e-3
rk3845 n949__vddio n38__vddio 104.4e-3
rk3846 n38__vddio n35__vddio 1.1705
rk3847 n35__vddio n950__vddio 196.8e-3
rk3848 n950__vddio n34__vddio 1.0796
rk3849 n34__vddio n951__vddio 437.6e-3
rk3850 n951__vddio n948__vddio 8.8496
rk3851 n758__vddio n31__vddio 441.3e-3
rk3852 n31__vddio n953__vddio 527.6e-3
rk3853 n953__vddio n30__vddio 111.9e-3
rk3854 n30__vddio n27__vddio 1.1771
rk3855 n27__vddio n954__vddio 200.1e-3
rk3856 n954__vddio n26__vddio 1.083
rk3857 n26__vddio n955__vddio 440.9e-3
rk3858 n955__vddio n952__vddio 8.8496
rk3859 n760__vddio n23__vddio 441.3e-3
rk3860 n23__vddio n957__vddio 527.6e-3
rk3861 n957__vddio n22__vddio 111.9e-3
rk3862 n22__vddio n19__vddio 1.1771
rk3863 n19__vddio n958__vddio 200.1e-3
rk3864 n958__vddio n18__vddio 1.083
rk3865 n18__vddio n959__vddio 440.9e-3
rk3866 n959__vddio n956__vddio 8.8496
rk3867 n761__vddio n15__vddio 444.1e-3
rk3868 n15__vddio n961__vddio 530.3e-3
rk3869 n961__vddio n14__vddio 116e-3
rk3870 n14__vddio n11__vddio 1.1827
rk3871 n11__vddio n962__vddio 202.9e-3
rk3872 n962__vddio n10__vddio 1.0857
rk3873 n10__vddio n963__vddio 443.7e-3
rk3874 n963__vddio n960__vddio 8.8496
rk3875 n686__vddio n687__vddio 7.5
rk3876 n686__vddio n689__vddio 3.75
rk3877 n686__vddio n690__vddio 3.75
rk3878 n686__vddio n691__vddio 3.75
rk3879 n686__vddio n692__vddio 3.75
rk3880 n686__vddio n693__vddio 3.75
rk3881 n686__vddio n694__vddio 3.75
rk3882 n686__vddio n695__vddio 3.75
rk3883 n686__vddio n696__vddio 3.75
rk3884 n686__vddio n697__vddio 3.75
rk3885 n699__vddio n700__vddio 3.1
rk3886 n686__vddio n704__vddio 3.75
rk3887 n686__vddio n708__vddio 3.75
rk3888 n686__vddio n712__vddio 3.75
rk3889 n686__vddio n716__vddio 3.75
rk3890 n686__vddio n720__vddio 3.75
rk3891 n686__vddio n725__vddio 3.75
rk3892 n686__vddio n729__vddio 3.75
rk3893 n686__vddio n734__vddio 3.75
rk3894 n686__vddio n738__vddio 3.75
rk3895 n686__vddio n742__vddio 3.75
rk3896 n686__vddio n746__vddio 3.75
rk3897 n686__vddio n750__vddio 3.75
rk3898 n686__vddio n755__vddio 3.75
rk3899 n686__vddio n759__vddio 3.75
rk3900 n762__vddio n763__vddio 3.1
rk3901 n762__vddio n764__vddio 3.1
rk3902 n762__vddio n765__vddio 3.1
rk3903 n699__vddio n766__vddio 3.1
rk3904 n699__vddio n767__vddio 3.1
rk3905 n768__vddio n769__vddio 3.1
rk3906 n768__vddio n770__vddio 3.1
rk3907 n768__vddio n771__vddio 3.1
rk3908 n772__vddio n773__vddio 3.1
rk3909 n772__vddio n774__vddio 3.1
rk3910 n772__vddio n775__vddio 3.1
rk3911 n776__vddio n777__vddio 3.1
rk3912 n776__vddio n778__vddio 3.1
rk3913 n776__vddio n779__vddio 3.1
rk3914 n780__vddio n781__vddio 3.1
rk3915 n780__vddio n782__vddio 3.1
rk3916 n780__vddio n783__vddio 3.1
rk3917 n784__vddio n785__vddio 3.1
rk3918 n784__vddio n786__vddio 3.1
rk3919 n784__vddio n787__vddio 3.1
rk3920 n788__vddio n789__vddio 3.1
rk3921 n788__vddio n790__vddio 3.1
rk3922 n788__vddio n791__vddio 3.1
rk3923 n792__vddio n793__vddio 3.1
rk3924 n792__vddio n794__vddio 3.1
rk3925 n792__vddio n795__vddio 3.1
rk3926 n796__vddio n797__vddio 3.1
rk3927 n796__vddio n798__vddio 3.1
rk3928 n796__vddio n799__vddio 3.1
rk3929 n800__vddio n801__vddio 3.1
rk3930 n800__vddio n802__vddio 3.1
rk3931 n800__vddio n803__vddio 3.1
rk3932 n804__vddio n805__vddio 3.1
rk3933 n804__vddio n806__vddio 3.1
rk3934 n804__vddio n807__vddio 3.1
rk3935 n808__vddio n809__vddio 3.1
rk3936 n808__vddio n810__vddio 3.1
rk3937 n808__vddio n811__vddio 3.1
rk3938 n812__vddio n813__vddio 3.1
rk3939 n812__vddio n814__vddio 3.1
rk3940 n812__vddio n815__vddio 3.1
rk3941 n816__vddio n817__vddio 3.1
rk3942 n816__vddio n818__vddio 3.1
rk3943 n816__vddio n819__vddio 3.1
rk3944 n820__vddio n821__vddio 3.1
rk3945 n820__vddio n822__vddio 3.1
rk3946 n820__vddio n823__vddio 3.1
rk3947 n824__vddio n825__vddio 3.1
rk3948 n824__vddio n826__vddio 3.1
rk3949 n824__vddio n827__vddio 3.1
rk3950 n828__vddio n829__vddio 3.1
rk3951 n828__vddio n830__vddio 3.1
rk3952 n828__vddio n831__vddio 3.1
rk3953 n832__vddio n833__vddio 3.1
rk3954 n832__vddio n834__vddio 3.1
rk3955 n832__vddio n835__vddio 3.1
rk3956 n836__vddio n837__vddio 3.1
rk3957 n836__vddio n838__vddio 3.1
rk3958 n836__vddio n839__vddio 3.1
rk3959 n840__vddio n841__vddio 3.1
rk3960 n840__vddio n842__vddio 3.1
rk3961 n840__vddio n843__vddio 3.1
rk3962 n844__vddio n845__vddio 3.1
rk3963 n844__vddio n846__vddio 3.1
rk3964 n844__vddio n847__vddio 3.1
rk3965 n848__vddio n849__vddio 3.1
rk3966 n848__vddio n850__vddio 3.1
rk3967 n848__vddio n851__vddio 3.1
rk3968 n852__vddio n853__vddio 3.1
rk3969 n852__vddio n854__vddio 3.1
rk3970 n852__vddio n855__vddio 3.1
rk3971 n856__vddio n857__vddio 3.1
rk3972 n856__vddio n858__vddio 3.1
rk3973 n856__vddio n859__vddio 3.1
rk3974 n860__vddio n861__vddio 3.1
rk3975 n860__vddio n862__vddio 3.1
rk3976 n860__vddio n863__vddio 3.1
rk3977 n864__vddio n865__vddio 3.1
rk3978 n864__vddio n866__vddio 3.1
rk3979 n864__vddio n867__vddio 3.1
rk3980 n868__vddio n869__vddio 3.1
rk3981 n868__vddio n870__vddio 3.1
rk3982 n868__vddio n871__vddio 3.1
rk3983 n872__vddio n873__vddio 3.1
rk3984 n872__vddio n874__vddio 3.1
rk3985 n872__vddio n875__vddio 3.1
rk3986 n876__vddio n877__vddio 3.1
rk3987 n876__vddio n878__vddio 3.1
rk3988 n876__vddio n879__vddio 3.1
rk3989 n880__vddio n881__vddio 3.1
rk3990 n880__vddio n882__vddio 3.1
rk3991 n880__vddio n883__vddio 3.1
rk3992 n884__vddio n885__vddio 3.1
rk3993 n884__vddio n886__vddio 3.1
rk3994 n884__vddio n887__vddio 3.1
rk3995 n888__vddio n889__vddio 3.1
rk3996 n888__vddio n890__vddio 3.1
rk3997 n888__vddio n891__vddio 3.1
rk3998 n892__vddio n893__vddio 3.1
rk3999 n892__vddio n894__vddio 3.1
rk4000 n892__vddio n895__vddio 3.1
rk4001 n896__vddio n897__vddio 3.1
rk4002 n896__vddio n898__vddio 3.1
rk4003 n896__vddio n899__vddio 3.1
rk4004 n900__vddio n901__vddio 3.1
rk4005 n900__vddio n902__vddio 3.1
rk4006 n900__vddio n903__vddio 3.1
rk4007 n904__vddio n905__vddio 3.1
rk4008 n904__vddio n906__vddio 3.1
rk4009 n904__vddio n907__vddio 3.1
rk4010 n908__vddio n909__vddio 3.1
rk4011 n908__vddio n910__vddio 3.1
rk4012 n908__vddio n911__vddio 3.1
rk4013 n912__vddio n913__vddio 3.1
rk4014 n912__vddio n914__vddio 3.1
rk4015 n912__vddio n915__vddio 3.1
rk4016 n916__vddio n917__vddio 3.1
rk4017 n916__vddio n918__vddio 3.1
rk4018 n916__vddio n919__vddio 3.1
rk4019 n920__vddio n921__vddio 3.1
rk4020 n920__vddio n922__vddio 3.1
rk4021 n920__vddio n923__vddio 3.1
rk4022 n924__vddio n925__vddio 3.1
rk4023 n924__vddio n926__vddio 3.1
rk4024 n924__vddio n927__vddio 3.1
rk4025 n928__vddio n929__vddio 3.1
rk4026 n928__vddio n930__vddio 3.1
rk4027 n928__vddio n931__vddio 3.1
rk4028 n932__vddio n933__vddio 3.1
rk4029 n932__vddio n934__vddio 3.1
rk4030 n932__vddio n935__vddio 3.1
rk4031 n936__vddio n937__vddio 3.1
rk4032 n936__vddio n938__vddio 3.1
rk4033 n936__vddio n939__vddio 3.1
rk4034 n940__vddio n941__vddio 3.1
rk4035 n940__vddio n942__vddio 3.1
rk4036 n940__vddio n943__vddio 3.1
rk4037 n944__vddio n945__vddio 3.1
rk4038 n944__vddio n946__vddio 3.1
rk4039 n944__vddio n947__vddio 3.1
rk4040 n948__vddio n949__vddio 3.1
rk4041 n948__vddio n950__vddio 3.1
rk4042 n948__vddio n951__vddio 3.1
rk4043 n952__vddio n953__vddio 3.1
rk4044 n952__vddio n954__vddio 3.1
rk4045 n952__vddio n955__vddio 3.1
rk4046 n956__vddio n957__vddio 3.1
rk4047 n956__vddio n958__vddio 3.1
rk4048 n956__vddio n959__vddio 3.1
rk4049 n960__vddio n961__vddio 3.1
rk4050 n960__vddio n962__vddio 3.1
rk4051 n960__vddio n963__vddio 3.1
rk4052 n1010__vss n1011__vss 37.6898
rk4053 n1011__vss n1012__vss 18.93e-3
rk4054 n1012__vss n1013__vss 105.1e-3
rk4055 n1013__vss n1014__vss 295.1e-3
rk4056 n1014__vss n1015__vss 173.2e-3
rk4057 n1011__vss n1016__vss 321.9e-3
rk4058 n1013__vss n1017__vss 75.1845
rk4059 n1014__vss n1018__vss 37.6898
rk4060 n1015__vss n1019__vss 37.6862
rk4061 n1015__vss n1020__vss 187.6e-3
rk4062 n1020__vss n1021__vss 37.6898
rk4063 n1020__vss n1022__vss 164.7e-3
rk4064 n1022__vss n1023__vss 37.6898
rk4065 n1022__vss n1024__vss 221.1e-3
rk4066 n1024__vss n1025__vss 260.6e-3
rk4067 n1025__vss n1026__vss 110.8e-3
rk4068 n1026__vss n1027__vss 202e-3
rk4069 n1027__vss n1028__vss 363.5e-3
rk4070 n1028__vss n1029__vss 126.4e-3
rk4071 n1029__vss n1030__vss 83.53e-3
rk4072 n1030__vss n1031__vss 76.35e-3
rk4073 n1031__vss n1032__vss 497.4e-3
rk4074 n1032__vss n1033__vss 18.93e-3
rk4075 n1033__vss n1034__vss 126.4e-3
rk4076 n1034__vss n1035__vss 159.9e-3
rk4077 n1035__vss n506__vss 88.67e-3
rk4078 n1025__vss n1036__vss 75.207
rk4079 n1026__vss n1037__vss 75.1361
rk4080 n1028__vss n1038__vss 75.207
rk4081 n1029__vss n1039__vss 75.212
rk4082 n1031__vss n1040__vss 37.6727
rk4083 n1033__vss n1041__vss 75.207
rk4084 n1034__vss n1042__vss 75.212
rk4085 n1035__vss n1043__vss 37.6727
rk4086 n506__vss n1044__vss 165.4e-3
rk4087 n1044__vss n1045__vss 248.6e-3
rk4088 n1045__vss n1046__vss 325.2e-3
rk4089 n1046__vss n1047__vss 191.2e-3
rk4090 n1047__vss n1048__vss 149.1e-3
rk4091 n1048__vss n1049__vss 110.8e-3
rk4092 n1049__vss n1050__vss 61.78e-3
rk4093 n1050__vss n1051__vss 59.6e-3
rk4094 n1051__vss n1052__vss 38.07e-3
rk4095 n1052__vss n1053__vss 79.72e-3
rk4096 n1053__vss n434__vss 57.94e-3
rk4097 n434__vss n1054__vss 170.4e-3
rk4098 n1054__vss n418__vss 354.6e-3
rk4099 n418__vss n1056__vss 235.4e-3
rk4100 n1056__vss n419__vss 274e-3
rk4101 n419__vss n1057__vss 858e-3
rk4102 n1057__vss n422__vss 78.33e-3
rk4103 n422__vss n423__vss 913.9e-3
rk4104 n423__vss n1055__vss 4.2519
rk4105 n1045__vss n1058__vss 75.207
rk4106 n1047__vss n1059__vss 75.207
rk4107 n1048__vss n1060__vss 37.6727
rk4108 n1049__vss n1061__vss 37.6727
rk4109 n1050__vss n1062__vss 37.6727
rk4110 n1052__vss n1063__vss 37.6727
rk4111 n1053__vss n1064__vss 75.2027
rk4112 n1054__vss n1065__vss 115.6e-3
rk4113 n1065__vss n1066__vss 48.62e-3
rk4114 n1066__vss n394__vss 351.3e-3
rk4115 n394__vss n1068__vss 232.1e-3
rk4116 n1068__vss n395__vss 270.6e-3
rk4117 n395__vss n1069__vss 856.6e-3
rk4118 n1069__vss n398__vss 73.07e-3
rk4119 n398__vss n399__vss 907.2e-3
rk4120 n399__vss n1067__vss 4.2486
rk4121 n1065__vss n1070__vss 37.6727
rk4122 n1066__vss n407__vss 26.1e-3
rk4123 n407__vss n1071__vss 32.3e-3
rk4124 n1071__vss n1072__vss 52.42e-3
rk4125 n1072__vss n1073__vss 55.8e-3
rk4126 n1073__vss n385__vss 351.3e-3
rk4127 n385__vss n1075__vss 232.1e-3
rk4128 n1075__vss n388__vss 270.6e-3
rk4129 n388__vss n1076__vss 856.6e-3
rk4130 n1076__vss n389__vss 73.07e-3
rk4131 n389__vss n392__vss 907.2e-3
rk4132 n392__vss n1074__vss 4.2486
rk4133 n1071__vss n1077__vss 37.6691
rk4134 n1072__vss n1078__vss 75.207
rk4135 n1073__vss n1079__vss 54.6e-3
rk4136 n1079__vss n1080__vss 112e-3
rk4137 n1080__vss n378__vss 354.6e-3
rk4138 n378__vss n1082__vss 235.4e-3
rk4139 n1082__vss n379__vss 274e-3
rk4140 n379__vss n1083__vss 858e-3
rk4141 n1083__vss n382__vss 78.33e-3
rk4142 n382__vss n383__vss 913.9e-3
rk4143 n383__vss n1081__vss 4.2519
rk4144 n1079__vss n1084__vss 75.2047
rk4145 n1080__vss n1085__vss 167.1e-3
rk4146 n1085__vss n370__vss 354.6e-3
rk4147 n370__vss n1087__vss 235.4e-3
rk4148 n1087__vss n371__vss 274e-3
rk4149 n371__vss n1088__vss 858e-3
rk4150 n1088__vss n374__vss 78.33e-3
rk4151 n374__vss n375__vss 913.9e-3
rk4152 n375__vss n1086__vss 4.2519
rk4153 n1085__vss n1089__vss 130.2e-3
rk4154 n1089__vss n1090__vss 36.87e-3
rk4155 n1090__vss n362__vss 354.6e-3
rk4156 n362__vss n1092__vss 235.4e-3
rk4157 n1092__vss n363__vss 274e-3
rk4158 n363__vss n1093__vss 858e-3
rk4159 n1093__vss n366__vss 78.33e-3
rk4160 n366__vss n367__vss 913.9e-3
rk4161 n367__vss n1091__vss 4.2519
rk4162 n1089__vss n1094__vss 37.6691
rk4163 n1090__vss n1095__vss 70.15e-3
rk4164 n1095__vss n1096__vss 61.78e-3
rk4165 n1096__vss n1097__vss 34.27e-3
rk4166 n1097__vss n354__vss 354.6e-3
rk4167 n354__vss n1099__vss 235.4e-3
rk4168 n1099__vss n355__vss 274e-3
rk4169 n355__vss n1100__vss 858e-3
rk4170 n1100__vss n358__vss 78.33e-3
rk4171 n358__vss n359__vss 913.9e-3
rk4172 n359__vss n1098__vss 4.2519
rk4173 n1095__vss n1101__vss 37.6727
rk4174 n1096__vss n1102__vss 37.6727
rk4175 n1097__vss n1103__vss 62.98e-3
rk4176 n1103__vss n1104__vss 79.72e-3
rk4177 n1104__vss n1105__vss 23.5e-3
rk4178 n1105__vss n345__vss 357.4e-3
rk4179 n345__vss n1107__vss 238.2e-3
rk4180 n1107__vss n348__vss 276.7e-3
rk4181 n348__vss n1108__vss 860.7e-3
rk4182 n1108__vss n349__vss 81.17e-3
rk4183 n349__vss n352__vss 919.4e-3
rk4184 n352__vss n1106__vss 4.2546
rk4185 n1103__vss n1109__vss 37.6727
rk4186 n1104__vss n1110__vss 75.2027
rk4187 n1105__vss n1111__vss 167.1e-3
rk4188 n1111__vss n338__vss 357.4e-3
rk4189 n338__vss n1113__vss 238.2e-3
rk4190 n1113__vss n339__vss 276.7e-3
rk4191 n339__vss n1114__vss 860.7e-3
rk4192 n1114__vss n342__vss 81.17e-3
rk4193 n342__vss n343__vss 919.4e-3
rk4194 n343__vss n1112__vss 4.2546
rk4195 n1111__vss n1115__vss 34.48e-3
rk4196 n1115__vss n1116__vss 121.8e-3
rk4197 n1116__vss n1117__vss 12.22e-3
rk4198 n1117__vss n330__vss 355.6e-3
rk4199 n330__vss n1119__vss 231.2e-3
rk4200 n1119__vss n331__vss 269.8e-3
rk4201 n331__vss n1120__vss 856.5e-3
rk4202 n1120__vss n334__vss 71.5e-3
rk4203 n334__vss n335__vss 905.5e-3
rk4204 n335__vss n1118__vss 4.2477
rk4205 n1116__vss n1121__vss 37.6727
rk4206 n1117__vss n1122__vss 85.2e-3
rk4207 n1122__vss n1123__vss 61.78e-3
rk4208 n1123__vss n1124__vss 17.52e-3
rk4209 n1124__vss n322__vss 350.5e-3
rk4210 n322__vss n1126__vss 231.2e-3
rk4211 n1126__vss n323__vss 269.8e-3
rk4212 n323__vss n1127__vss 856.5e-3
rk4213 n1127__vss n326__vss 71.5e-3
rk4214 n326__vss n327__vss 905.5e-3
rk4215 n327__vss n1125__vss 4.2477
rk4216 n1122__vss n1128__vss 37.6727
rk4217 n1123__vss n1129__vss 75.207
rk4218 n1124__vss n1130__vss 92.88e-3
rk4219 n1130__vss n1131__vss 73.74e-3
rk4220 n1131__vss n314__vss 357.4e-3
rk4221 n314__vss n1133__vss 238.2e-3
rk4222 n1133__vss n315__vss 276.7e-3
rk4223 n315__vss n1134__vss 860.7e-3
rk4224 n1134__vss n318__vss 81.17e-3
rk4225 n318__vss n319__vss 919.4e-3
rk4226 n319__vss n1132__vss 4.2546
rk4227 n1130__vss n1135__vss 75.2047
rk4228 n1131__vss n1136__vss 106.3e-3
rk4229 n1136__vss n1137__vss 60.8e-3
rk4230 n1137__vss n306__vss 357.4e-3
rk4231 n306__vss n1139__vss 238.2e-3
rk4232 n1139__vss n307__vss 276.7e-3
rk4233 n307__vss n1140__vss 860.7e-3
rk4234 n1140__vss n310__vss 81.17e-3
rk4235 n310__vss n311__vss 919.4e-3
rk4236 n311__vss n1138__vss 4.2546
rk4237 n1137__vss n1141__vss 167.1e-3
rk4238 n1141__vss n298__vss 354.6e-3
rk4239 n298__vss n1143__vss 235.4e-3
rk4240 n1143__vss n299__vss 274e-3
rk4241 n299__vss n1144__vss 858e-3
rk4242 n1144__vss n302__vss 78.33e-3
rk4243 n302__vss n303__vss 913.9e-3
rk4244 n303__vss n1142__vss 4.2519
rk4245 n1141__vss n1145__vss 167.1e-3
rk4246 n1145__vss n290__vss 354.6e-3
rk4247 n290__vss n1147__vss 235.4e-3
rk4248 n1147__vss n291__vss 274e-3
rk4249 n291__vss n1148__vss 858e-3
rk4250 n1148__vss n294__vss 78.33e-3
rk4251 n294__vss n295__vss 913.9e-3
rk4252 n295__vss n1146__vss 4.2519
rk4253 n1145__vss n1149__vss 178e-3
rk4254 n1149__vss n282__vss 353.8e-3
rk4255 n282__vss n1151__vss 238.2e-3
rk4256 n1151__vss n283__vss 276.7e-3
rk4257 n283__vss n1152__vss 860.7e-3
rk4258 n1152__vss n286__vss 81.17e-3
rk4259 n286__vss n287__vss 919.4e-3
rk4260 n287__vss n1150__vss 4.2546
rk4261 n1149__vss n1153__vss 156.5e-3
rk4262 n1153__vss n274__vss 357.4e-3
rk4263 n274__vss n1155__vss 238.2e-3
rk4264 n1155__vss n275__vss 276.7e-3
rk4265 n275__vss n1156__vss 860.7e-3
rk4266 n1156__vss n278__vss 81.17e-3
rk4267 n278__vss n279__vss 919.4e-3
rk4268 n279__vss n1154__vss 4.2546
rk4269 n1153__vss n1157__vss 167.1e-3
rk4270 n1157__vss n266__vss 350.5e-3
rk4271 n266__vss n1159__vss 231.2e-3
rk4272 n1159__vss n267__vss 269.8e-3
rk4273 n267__vss n1160__vss 856.5e-3
rk4274 n1160__vss n270__vss 71.5e-3
rk4275 n270__vss n271__vss 905.5e-3
rk4276 n271__vss n1158__vss 4.2477
rk4277 n1157__vss n1161__vss 167.1e-3
rk4278 n1161__vss n258__vss 350.5e-3
rk4279 n258__vss n1163__vss 231.2e-3
rk4280 n1163__vss n259__vss 269.8e-3
rk4281 n259__vss n1164__vss 856.5e-3
rk4282 n1164__vss n262__vss 71.5e-3
rk4283 n262__vss n263__vss 905.5e-3
rk4284 n263__vss n1162__vss 4.2477
rk4285 n1161__vss n1165__vss 82.33e-3
rk4286 n1165__vss n1166__vss 84.72e-3
rk4287 n1166__vss n250__vss 357.4e-3
rk4288 n250__vss n1168__vss 238.2e-3
rk4289 n1168__vss n251__vss 276.7e-3
rk4290 n251__vss n1169__vss 860.7e-3
rk4291 n1169__vss n254__vss 81.17e-3
rk4292 n254__vss n255__vss 919.4e-3
rk4293 n255__vss n1167__vss 4.2546
rk4294 n1166__vss n1170__vss 167.1e-3
rk4295 n1170__vss n242__vss 354.6e-3
rk4296 n242__vss n1172__vss 235.4e-3
rk4297 n1172__vss n243__vss 274e-3
rk4298 n243__vss n1173__vss 858e-3
rk4299 n1173__vss n246__vss 78.33e-3
rk4300 n246__vss n247__vss 913.9e-3
rk4301 n247__vss n1171__vss 4.2519
rk4302 n1170__vss n1174__vss 167.1e-3
rk4303 n1174__vss n234__vss 354.6e-3
rk4304 n234__vss n1176__vss 235.4e-3
rk4305 n1176__vss n235__vss 274e-3
rk4306 n235__vss n1177__vss 858e-3
rk4307 n1177__vss n238__vss 78.33e-3
rk4308 n238__vss n239__vss 913.9e-3
rk4309 n239__vss n1175__vss 4.2519
rk4310 n1174__vss n1178__vss 154.1e-3
rk4311 n1178__vss n226__vss 353.8e-3
rk4312 n226__vss n1180__vss 238.2e-3
rk4313 n1180__vss n227__vss 276.7e-3
rk4314 n227__vss n1181__vss 860.7e-3
rk4315 n1181__vss n230__vss 81.17e-3
rk4316 n230__vss n231__vss 919.4e-3
rk4317 n231__vss n1179__vss 4.2546
rk4318 n1178__vss n1182__vss 180.4e-3
rk4319 n1182__vss n218__vss 357.4e-3
rk4320 n218__vss n1184__vss 238.2e-3
rk4321 n1184__vss n219__vss 276.7e-3
rk4322 n219__vss n1185__vss 860.7e-3
rk4323 n1185__vss n222__vss 81.17e-3
rk4324 n222__vss n223__vss 919.4e-3
rk4325 n223__vss n1183__vss 4.2546
rk4326 n1182__vss n1186__vss 167.1e-3
rk4327 n1186__vss n210__vss 350.5e-3
rk4328 n210__vss n1188__vss 231.2e-3
rk4329 n1188__vss n211__vss 269.8e-3
rk4330 n211__vss n1189__vss 856.5e-3
rk4331 n1189__vss n214__vss 71.5e-3
rk4332 n214__vss n215__vss 905.5e-3
rk4333 n215__vss n1187__vss 4.2477
rk4334 n1186__vss n1190__vss 167.1e-3
rk4335 n1190__vss n202__vss 350.5e-3
rk4336 n202__vss n1192__vss 231.2e-3
rk4337 n1192__vss n203__vss 269.8e-3
rk4338 n203__vss n1193__vss 856.5e-3
rk4339 n1193__vss n206__vss 71.5e-3
rk4340 n206__vss n207__vss 905.5e-3
rk4341 n207__vss n1191__vss 4.2477
rk4342 n1190__vss n1194__vss 58.4e-3
rk4343 n1194__vss n1195__vss 108.6e-3
rk4344 n1195__vss n194__vss 357.4e-3
rk4345 n194__vss n1197__vss 238.2e-3
rk4346 n1197__vss n195__vss 276.7e-3
rk4347 n195__vss n1198__vss 860.7e-3
rk4348 n1198__vss n198__vss 81.17e-3
rk4349 n198__vss n199__vss 919.4e-3
rk4350 n199__vss n1196__vss 4.2546
rk4351 n1195__vss n1199__vss 167.1e-3
rk4352 n1199__vss n186__vss 357.4e-3
rk4353 n186__vss n1201__vss 238.2e-3
rk4354 n1201__vss n187__vss 276.7e-3
rk4355 n187__vss n1202__vss 860.7e-3
rk4356 n1202__vss n190__vss 81.17e-3
rk4357 n190__vss n191__vss 919.4e-3
rk4358 n191__vss n1200__vss 4.2546
rk4359 n1199__vss n1203__vss 167.1e-3
rk4360 n1203__vss n178__vss 354.6e-3
rk4361 n178__vss n1205__vss 235.4e-3
rk4362 n1205__vss n179__vss 274e-3
rk4363 n179__vss n1206__vss 858e-3
rk4364 n1206__vss n182__vss 78.33e-3
rk4365 n182__vss n183__vss 913.9e-3
rk4366 n183__vss n1204__vss 4.2519
rk4367 n1203__vss n1207__vss 130.2e-3
rk4368 n1207__vss n1208__vss 36.87e-3
rk4369 n1208__vss n170__vss 354.6e-3
rk4370 n170__vss n1210__vss 235.4e-3
rk4371 n1210__vss n171__vss 274e-3
rk4372 n171__vss n1211__vss 858e-3
rk4373 n1211__vss n174__vss 78.33e-3
rk4374 n174__vss n175__vss 913.9e-3
rk4375 n175__vss n1209__vss 4.2519
rk4376 n1208__vss n1212__vss 167.1e-3
rk4377 n1212__vss n162__vss 357.4e-3
rk4378 n162__vss n1214__vss 238.2e-3
rk4379 n1214__vss n163__vss 276.7e-3
rk4380 n163__vss n1215__vss 860.7e-3
rk4381 n1215__vss n166__vss 81.17e-3
rk4382 n166__vss n167__vss 919.4e-3
rk4383 n167__vss n1213__vss 4.2546
rk4384 n1212__vss n1216__vss 167.1e-3
rk4385 n1216__vss n154__vss 357.4e-3
rk4386 n154__vss n1218__vss 238.2e-3
rk4387 n1218__vss n155__vss 276.7e-3
rk4388 n155__vss n1219__vss 860.7e-3
rk4389 n1219__vss n158__vss 81.17e-3
rk4390 n158__vss n159__vss 919.4e-3
rk4391 n159__vss n1217__vss 4.2546
rk4392 n1216__vss n1220__vss 167.1e-3
rk4393 n1220__vss n146__vss 350.5e-3
rk4394 n146__vss n1222__vss 231.2e-3
rk4395 n1222__vss n147__vss 269.8e-3
rk4396 n147__vss n1223__vss 856.5e-3
rk4397 n1223__vss n150__vss 71.5e-3
rk4398 n150__vss n151__vss 905.5e-3
rk4399 n151__vss n1221__vss 4.2477
rk4400 n1220__vss n1224__vss 34.48e-3
rk4401 n1224__vss n1225__vss 132.6e-3
rk4402 n1225__vss n138__vss 350.5e-3
rk4403 n138__vss n1227__vss 231.2e-3
rk4404 n1227__vss n139__vss 269.8e-3
rk4405 n139__vss n1228__vss 856.5e-3
rk4406 n1228__vss n142__vss 71.5e-3
rk4407 n142__vss n143__vss 905.5e-3
rk4408 n143__vss n1226__vss 4.2477
rk4409 n1225__vss n1229__vss 167.1e-3
rk4410 n1229__vss n130__vss 357.4e-3
rk4411 n130__vss n1231__vss 238.2e-3
rk4412 n1231__vss n131__vss 276.7e-3
rk4413 n131__vss n1232__vss 860.7e-3
rk4414 n1232__vss n134__vss 81.17e-3
rk4415 n134__vss n135__vss 919.4e-3
rk4416 n135__vss n1230__vss 4.2546
rk4417 n1229__vss n1233__vss 167.1e-3
rk4418 n1233__vss n122__vss 355.5e-3
rk4419 n122__vss n1235__vss 236.3e-3
rk4420 n1235__vss n123__vss 274.8e-3
rk4421 n123__vss n1236__vss 857e-3
rk4422 n1236__vss n126__vss 81.17e-3
rk4423 n126__vss n127__vss 915.7e-3
rk4424 n127__vss n1234__vss 4.2528
rk4425 n1233__vss n1237__vss 106.3e-3
rk4426 n1237__vss n1238__vss 60.8e-3
rk4427 n1238__vss n114__vss 355.5e-3
rk4428 n114__vss n1240__vss 236.3e-3
rk4429 n1240__vss n115__vss 274.8e-3
rk4430 n115__vss n1241__vss 857e-3
rk4431 n1241__vss n118__vss 81.17e-3
rk4432 n118__vss n119__vss 915.7e-3
rk4433 n119__vss n1239__vss 4.2528
rk4434 n1238__vss n1242__vss 167.1e-3
rk4435 n1242__vss n106__vss 351.3e-3
rk4436 n106__vss n1244__vss 232.1e-3
rk4437 n1244__vss n107__vss 270.6e-3
rk4438 n107__vss n1245__vss 856.6e-3
rk4439 n1245__vss n110__vss 73.07e-3
rk4440 n110__vss n111__vss 907.2e-3
rk4441 n111__vss n1243__vss 4.2486
rk4442 n1242__vss n1246__vss 167.1e-3
rk4443 n1246__vss n98__vss 351.3e-3
rk4444 n98__vss n1248__vss 232.1e-3
rk4445 n1248__vss n99__vss 270.6e-3
rk4446 n99__vss n1249__vss 856.6e-3
rk4447 n1249__vss n102__vss 73.07e-3
rk4448 n102__vss n103__vss 907.2e-3
rk4449 n103__vss n1247__vss 4.2486
rk4450 n1246__vss n1250__vss 178e-3
rk4451 n1250__vss n90__vss 351e-3
rk4452 n90__vss n1252__vss 235.4e-3
rk4453 n1252__vss n91__vss 274e-3
rk4454 n91__vss n1253__vss 858e-3
rk4455 n1253__vss n94__vss 78.33e-3
rk4456 n94__vss n95__vss 913.9e-3
rk4457 n95__vss n1251__vss 4.2519
rk4458 n1250__vss n1254__vss 156.5e-3
rk4459 n1254__vss n82__vss 354.6e-3
rk4460 n82__vss n1256__vss 235.4e-3
rk4461 n1256__vss n83__vss 274e-3
rk4462 n83__vss n1257__vss 858e-3
rk4463 n1257__vss n86__vss 78.33e-3
rk4464 n86__vss n87__vss 913.9e-3
rk4465 n87__vss n1255__vss 4.2519
rk4466 n1254__vss n1258__vss 167.1e-3
rk4467 n1258__vss n74__vss 357.4e-3
rk4468 n74__vss n1260__vss 238.2e-3
rk4469 n1260__vss n75__vss 276.7e-3
rk4470 n75__vss n1261__vss 860.7e-3
rk4471 n1261__vss n78__vss 81.17e-3
rk4472 n78__vss n79__vss 919.4e-3
rk4473 n79__vss n1259__vss 4.2546
rk4474 n1258__vss n1262__vss 167.1e-3
rk4475 n1262__vss n66__vss 357.4e-3
rk4476 n66__vss n1264__vss 238.2e-3
rk4477 n1264__vss n67__vss 276.7e-3
rk4478 n67__vss n1265__vss 860.7e-3
rk4479 n1265__vss n70__vss 81.17e-3
rk4480 n70__vss n71__vss 919.4e-3
rk4481 n71__vss n1263__vss 4.2546
rk4482 n1262__vss n1266__vss 82.33e-3
rk4483 n1266__vss n1267__vss 84.72e-3
rk4484 n1267__vss n58__vss 355.5e-3
rk4485 n58__vss n1269__vss 236.3e-3
rk4486 n1269__vss n59__vss 274.8e-3
rk4487 n59__vss n1270__vss 857e-3
rk4488 n1270__vss n62__vss 81.17e-3
rk4489 n62__vss n63__vss 915.7e-3
rk4490 n63__vss n1268__vss 4.2528
rk4491 n1267__vss n1271__vss 167.1e-3
rk4492 n1271__vss n50__vss 355.5e-3
rk4493 n50__vss n1273__vss 236.3e-3
rk4494 n1273__vss n51__vss 274.8e-3
rk4495 n51__vss n1274__vss 857e-3
rk4496 n1274__vss n54__vss 81.17e-3
rk4497 n54__vss n55__vss 915.7e-3
rk4498 n55__vss n1272__vss 4.2528
rk4499 n1271__vss n1275__vss 167.1e-3
rk4500 n1275__vss n42__vss 351.3e-3
rk4501 n42__vss n1277__vss 232.1e-3
rk4502 n1277__vss n43__vss 270.6e-3
rk4503 n43__vss n1278__vss 856.6e-3
rk4504 n1278__vss n46__vss 73.07e-3
rk4505 n46__vss n47__vss 907.2e-3
rk4506 n47__vss n1276__vss 4.2486
rk4507 n1275__vss n1279__vss 154.1e-3
rk4508 n1279__vss n34__vss 347.7e-3
rk4509 n34__vss n1281__vss 232.1e-3
rk4510 n1281__vss n35__vss 270.6e-3
rk4511 n35__vss n1282__vss 856.6e-3
rk4512 n1282__vss n38__vss 73.07e-3
rk4513 n38__vss n39__vss 907.2e-3
rk4514 n39__vss n1280__vss 4.2486
rk4515 n1279__vss n1283__vss 180.4e-3
rk4516 n1283__vss n26__vss 354.6e-3
rk4517 n26__vss n1285__vss 235.4e-3
rk4518 n1285__vss n27__vss 274e-3
rk4519 n27__vss n1286__vss 858e-3
rk4520 n1286__vss n30__vss 78.33e-3
rk4521 n30__vss n31__vss 913.9e-3
rk4522 n31__vss n1284__vss 4.2519
rk4523 n1283__vss n1287__vss 167.1e-3
rk4524 n1287__vss n18__vss 354.6e-3
rk4525 n18__vss n1289__vss 235.4e-3
rk4526 n1289__vss n19__vss 274e-3
rk4527 n19__vss n1290__vss 858e-3
rk4528 n1290__vss n22__vss 78.33e-3
rk4529 n22__vss n23__vss 913.9e-3
rk4530 n23__vss n1288__vss 4.2519
rk4531 n1287__vss n1291__vss 167.1e-3
rk4532 n1291__vss n10__vss 357.4e-3
rk4533 n10__vss n1293__vss 238.2e-3
rk4534 n1293__vss n11__vss 276.7e-3
rk4535 n11__vss n1294__vss 860.7e-3
rk4536 n1294__vss n14__vss 81.17e-3
rk4537 n14__vss n15__vss 919.4e-3
rk4538 n15__vss n1292__vss 4.2546
rk4539 n1291__vss n2__vss 512.3e-3
rk4540 n2__vss n1296__vss 236.3e-3
rk4541 n1296__vss n3__vss 274.8e-3
rk4542 n3__vss n1297__vss 857e-3
rk4543 n1297__vss n6__vss 81.17e-3
rk4544 n6__vss n7__vss 915.7e-3
rk4545 n7__vss n1295__vss 4.2528
rk4546 n640__vss n1012__vss 3.1
rk4547 n640__vss n1015__vss 3.1
rk4548 n640__vss n1024__vss 3.1
rk4549 n640__vss n1027__vss 3.1
rk4550 n640__vss n1030__vss 3.1
rk4551 n640__vss n1032__vss 3.1
rk4552 n640__vss n1044__vss 3.1
rk4553 n640__vss n1046__vss 3.1
rk4554 n640__vss n1051__vss 3.1
rk4555 n1055__vss n1056__vss 7.5
rk4556 n1055__vss n1057__vss 3.75
rk4557 n1067__vss n1068__vss 7.5
rk4558 n1067__vss n1069__vss 3.75
rk4559 n640__vss n1071__vss 3.1
rk4560 n1074__vss n1075__vss 7.5
rk4561 n1074__vss n1076__vss 3.75
rk4562 n1081__vss n1082__vss 7.5
rk4563 n1081__vss n1083__vss 3.75
rk4564 n1086__vss n1087__vss 7.5
rk4565 n1086__vss n1088__vss 3.75
rk4566 n640__vss n1089__vss 3.1
rk4567 n1091__vss n1092__vss 7.5
rk4568 n1091__vss n1093__vss 3.75
rk4569 n1098__vss n1099__vss 7.5
rk4570 n1098__vss n1100__vss 3.75
rk4571 n1106__vss n1107__vss 7.5
rk4572 n1106__vss n1108__vss 3.75
rk4573 n1112__vss n1113__vss 7.5
rk4574 n1112__vss n1114__vss 3.75
rk4575 n640__vss n1115__vss 3.1
rk4576 n1118__vss n1119__vss 7.5
rk4577 n1118__vss n1120__vss 3.75
rk4578 n1125__vss n1126__vss 7.5
rk4579 n1125__vss n1127__vss 3.75
rk4580 n1132__vss n1133__vss 7.5
rk4581 n1132__vss n1134__vss 3.75
rk4582 n640__vss n1136__vss 3.1
rk4583 n1138__vss n1139__vss 7.5
rk4584 n1138__vss n1140__vss 3.75
rk4585 n1142__vss n1143__vss 7.5
rk4586 n1142__vss n1144__vss 3.75
rk4587 n1146__vss n1147__vss 7.5
rk4588 n1146__vss n1148__vss 3.75
rk4589 n640__vss n1149__vss 3.1
rk4590 n1150__vss n1151__vss 7.5
rk4591 n1150__vss n1152__vss 3.75
rk4592 n1154__vss n1155__vss 7.5
rk4593 n1154__vss n1156__vss 3.75
rk4594 n1158__vss n1159__vss 7.5
rk4595 n1158__vss n1160__vss 3.75
rk4596 n1162__vss n1163__vss 7.5
rk4597 n1162__vss n1164__vss 3.75
rk4598 n640__vss n1165__vss 3.1
rk4599 n1167__vss n1168__vss 7.5
rk4600 n1167__vss n1169__vss 3.75
rk4601 n1171__vss n1172__vss 7.5
rk4602 n1171__vss n1173__vss 3.75
rk4603 n1175__vss n1176__vss 7.5
rk4604 n1175__vss n1177__vss 3.75
rk4605 n640__vss n1178__vss 3.1
rk4606 n1179__vss n1180__vss 7.5
rk4607 n1179__vss n1181__vss 3.75
rk4608 n1183__vss n1184__vss 7.5
rk4609 n1183__vss n1185__vss 3.75
rk4610 n1187__vss n1188__vss 7.5
rk4611 n1187__vss n1189__vss 3.75
rk4612 n1191__vss n1192__vss 7.5
rk4613 n1191__vss n1193__vss 3.75
rk4614 n640__vss n1194__vss 3.1
rk4615 n1196__vss n1197__vss 7.5
rk4616 n1196__vss n1198__vss 3.75
rk4617 n1200__vss n1201__vss 7.5
rk4618 n1200__vss n1202__vss 3.75
rk4619 n1204__vss n1205__vss 7.5
rk4620 n1204__vss n1206__vss 3.75
rk4621 n640__vss n1207__vss 3.1
rk4622 n1209__vss n1210__vss 7.5
rk4623 n1209__vss n1211__vss 3.75
rk4624 n1213__vss n1214__vss 7.5
rk4625 n1213__vss n1215__vss 3.75
rk4626 n1217__vss n1218__vss 7.5
rk4627 n1217__vss n1219__vss 3.75
rk4628 n1221__vss n1222__vss 7.5
rk4629 n1221__vss n1223__vss 3.75
rk4630 n640__vss n1224__vss 3.1
rk4631 n1226__vss n1227__vss 7.5
rk4632 n1226__vss n1228__vss 3.75
rk4633 n1230__vss n1231__vss 7.5
rk4634 n1230__vss n1232__vss 3.75
rk4635 n1234__vss n1235__vss 7.5
rk4636 n1234__vss n1236__vss 3.75
rk4637 n640__vss n1237__vss 3.1
rk4638 n1239__vss n1240__vss 7.5
rk4639 n1239__vss n1241__vss 3.75
rk4640 n1243__vss n1244__vss 7.5
rk4641 n1243__vss n1245__vss 3.75
rk4642 n1247__vss n1248__vss 7.5
rk4643 n1247__vss n1249__vss 3.75
rk4644 n640__vss n1250__vss 3.1
rk4645 n1251__vss n1252__vss 7.5
rk4646 n1251__vss n1253__vss 3.75
rk4647 n1255__vss n1256__vss 7.5
rk4648 n1255__vss n1257__vss 3.75
rk4649 n1259__vss n1260__vss 7.5
rk4650 n1259__vss n1261__vss 3.75
rk4651 n1263__vss n1264__vss 7.5
rk4652 n1263__vss n1265__vss 3.75
rk4653 n640__vss n1266__vss 3.1
rk4654 n1268__vss n1269__vss 7.5
rk4655 n1268__vss n1270__vss 3.75
rk4656 n1272__vss n1273__vss 7.5
rk4657 n1272__vss n1274__vss 3.75
rk4658 n1276__vss n1277__vss 7.5
rk4659 n1276__vss n1278__vss 3.75
rk4660 n640__vss n1279__vss 3.1
rk4661 n1280__vss n1281__vss 7.5
rk4662 n1280__vss n1282__vss 3.75
rk4663 n1284__vss n1285__vss 7.5
rk4664 n1284__vss n1286__vss 3.75
rk4665 n1288__vss n1289__vss 7.5
rk4666 n1288__vss n1290__vss 3.75
rk4667 n1292__vss n1293__vss 7.5
rk4668 n1292__vss n1294__vss 3.75
rk4669 n1295__vss n1296__vss 7.5
rk4670 n1295__vss n1297__vss 3.75
rl1 i18__net5 n2__i18__net5 26.7741
rl2 n2__i18__net5 n3__i18__net5 29.8991
rl3 n4__i18__net5 n5__i18__net5 26.7741
rl4 n5__i18__net5 n6__i18__net5 29.8991
rl5 n7__i18__net5 n8__i18__net5 26.7741
rl6 n8__i18__net5 n9__i18__net5 29.8991
rl7 n10__i18__net5 n11__i18__net5 26.7741
rl8 n11__i18__net5 n12__i18__net5 29.8991
rl9 n13__i18__net5 n14__i18__net5 26.7741
rl10 n14__i18__net5 n15__i18__net5 29.8991
rl11 n16__i18__net5 n17__i18__net5 26.7741
rl12 n17__i18__net5 n18__i18__net5 29.8991
rl13 n19__i18__net5 n20__i18__net5 26.7741
rl14 n20__i18__net5 n21__i18__net5 29.8991
rl15 n22__i18__net5 n23__i18__net5 26.7741
rl16 n23__i18__net5 n24__i18__net5 29.8991
rl17 n25__i18__net5 n26__i18__net5 26.7741
rl18 n26__i18__net5 n27__i18__net5 29.8991
rl19 n28__i18__net5 n29__i18__net5 26.7741
rl20 n29__i18__net5 n30__i18__net5 29.8991
rl21 n31__i18__net5 n32__i18__net5 26.7741
rl22 n32__i18__net5 n33__i18__net5 29.8991
rl23 n34__i18__net5 n35__i18__net5 26.7741
rl24 n35__i18__net5 n36__i18__net5 29.8991
rl25 n37__i18__net5 n38__i18__net5 26.7741
rl26 n38__i18__net5 n39__i18__net5 29.8991
rl27 n40__i18__net5 n41__i18__net5 26.7741
rl28 n41__i18__net5 n42__i18__net5 29.8991
rl29 n43__i18__net5 n44__i18__net5 26.7741
rl30 n44__i18__net5 n45__i18__net5 29.8991
rl31 n50__i18__net5 n51__i18__net5 26.7741
rl32 n51__i18__net5 n52__i18__net5 29.8991
rl33 n53__i18__net5 n54__i18__net5 26.7741
rl34 n54__i18__net5 n55__i18__net5 29.8991
rl35 n60__i18__net5 n61__i18__net5 26.7741
rl36 n61__i18__net5 n62__i18__net5 29.8991
rl37 n63__i18__net5 n64__i18__net5 26.7741
rl38 n64__i18__net5 n65__i18__net5 29.8991
rl39 n68__i18__net5 n69__i18__net5 26.7741
rl40 n69__i18__net5 n70__i18__net5 29.8991
rl41 n73__i18__net5 n74__i18__net5 26.7741
rl42 n74__i18__net5 n75__i18__net5 29.8991
rl43 n78__i18__net5 n79__i18__net5 26.7741
rl44 n79__i18__net5 n80__i18__net5 29.8991
rl45 n85__i18__net5 n86__i18__net5 26.7741
rl46 n86__i18__net5 n87__i18__net5 29.8991
rl47 n90__i18__net5 n91__i18__net5 26.7741
rl48 n91__i18__net5 n92__i18__net5 29.8991
rl49 n95__i18__net5 n96__i18__net5 26.7741
rl50 n96__i18__net5 n97__i18__net5 29.8991
rl51 n100__i18__net5 n101__i18__net5 26.7741
rl52 n101__i18__net5 n102__i18__net5 29.8991
rl53 n103__i18__net5 n104__i18__net5 26.7741
rl54 n104__i18__net5 n105__i18__net5 29.8991
rl55 n110__i18__net5 n111__i18__net5 26.7741
rl56 n111__i18__net5 n112__i18__net5 29.8991
rl57 n115__i18__net5 n116__i18__net5 26.7741
rl58 n116__i18__net5 n117__i18__net5 29.8991
rl59 n120__i18__net5 n121__i18__net5 26.7741
rl60 n121__i18__net5 n122__i18__net5 29.8991
rl61 n123__i18__net5 n124__i18__net5 26.7741
rl62 n124__i18__net5 n125__i18__net5 29.8991
rl63 n129__i18__net5 n130__i18__net5 26.7741
rl64 n130__i18__net5 n131__i18__net5 29.8991
rl65 n135__i18__net5 n136__i18__net5 26.7741
rl66 n136__i18__net5 n137__i18__net5 29.8991
rl67 n138__i18__net5 n139__i18__net5 26.7741
rl68 n139__i18__net5 n140__i18__net5 29.8991
rl69 n143__i18__net5 n144__i18__net5 26.7741
rl70 n144__i18__net5 n145__i18__net5 29.8991
rl71 n148__i18__net5 n149__i18__net5 26.7741
rl72 n149__i18__net5 n150__i18__net5 29.8991
rl73 n153__i18__net5 n154__i18__net5 26.7741
rl74 n154__i18__net5 n155__i18__net5 29.8991
rl75 n160__i18__net5 n161__i18__net5 26.7741
rl76 n161__i18__net5 n162__i18__net5 29.8991
rl77 n164__i18__net5 n165__i18__net5 26.7741
rl78 n165__i18__net5 n166__i18__net5 29.8991
rl79 n170__i18__net5 n171__i18__net5 26.7741
rl80 n171__i18__net5 n172__i18__net5 29.8991
rl81 n173__i18__net5 n174__i18__net5 26.7741
rl82 n174__i18__net5 n175__i18__net5 29.8991
rl83 n179__i18__net5 n180__i18__net5 26.7741
rl84 n180__i18__net5 n181__i18__net5 29.8991
rl85 n185__i18__net5 n186__i18__net5 26.7741
rl86 n186__i18__net5 n187__i18__net5 29.8991
rl87 n188__i18__net5 n189__i18__net5 26.7741
rl88 n189__i18__net5 n190__i18__net5 29.8991
rl89 n193__i18__net5 n194__i18__net5 26.7741
rl90 n194__i18__net5 n195__i18__net5 29.8991
rl91 n199__i18__net5 n200__i18__net5 26.7741
rl92 n200__i18__net5 n201__i18__net5 29.8991
rl93 n203__i18__net5 n204__i18__net5 26.7741
rl94 n204__i18__net5 n205__i18__net5 29.8991
rl95 n208__i18__net5 n209__i18__net5 26.7741
rl96 n209__i18__net5 n210__i18__net5 29.8991
rl97 n214__i18__net5 n215__i18__net5 26.7741
rl98 n215__i18__net5 n216__i18__net5 29.8991
rl99 n218__i18__net5 n219__i18__net5 26.7741
rl100 n219__i18__net5 n220__i18__net5 29.8991
rl101 n223__i18__net5 n224__i18__net5 26.7741
rl102 n224__i18__net5 n225__i18__net5 29.8991
rl103 n228__i18__net5 n229__i18__net5 26.7741
rl104 n229__i18__net5 n230__i18__net5 29.8991
rl105 n235__i18__net5 n236__i18__net5 26.7741
rl106 n236__i18__net5 n237__i18__net5 29.8991
rl107 n240__i18__net5 n241__i18__net5 26.7741
rl108 n241__i18__net5 n242__i18__net5 29.8991
rl109 n245__i18__net5 n246__i18__net5 26.7741
rl110 n246__i18__net5 n247__i18__net5 29.8991
rl111 n250__i18__net5 n251__i18__net5 26.7741
rl112 n251__i18__net5 n252__i18__net5 29.8991
rl113 n253__i18__net5 n254__i18__net5 26.7741
rl114 n254__i18__net5 n255__i18__net5 29.8991
rl115 n258__i18__net5 n259__i18__net5 26.7741
rl116 n259__i18__net5 n260__i18__net5 29.8991
rl117 n265__i18__net5 n266__i18__net5 26.7741
rl118 n266__i18__net5 n267__i18__net5 29.8991
rl119 n268__i18__net5 n269__i18__net5 26.7741
rl120 n269__i18__net5 n270__i18__net5 29.8991
rl121 n275__i18__net5 n276__i18__net5 26.7741
rl122 n276__i18__net5 n277__i18__net5 29.8991
rl123 n278__i18__net5 n279__i18__net5 26.7741
rl124 n279__i18__net5 n280__i18__net5 29.8991
rl125 n283__i18__net5 n284__i18__net5 26.7741
rl126 n284__i18__net5 n285__i18__net5 29.8991
rl127 n288__i18__net5 n289__i18__net5 26.7741
rl128 n289__i18__net5 n290__i18__net5 29.8991
rl129 n293__i18__net5 n294__i18__net5 26.7741
rl130 n294__i18__net5 n295__i18__net5 29.8991
rl131 n298__i18__net5 n299__i18__net5 26.7741
rl132 n299__i18__net5 n300__i18__net5 29.8991
rl133 n303__i18__net5 n304__i18__net5 26.7741
rl134 n304__i18__net5 n305__i18__net5 29.8991
rl135 n310__i18__net5 n311__i18__net5 26.7741
rl136 n311__i18__net5 n312__i18__net5 29.8991
rl137 n313__i18__net5 n314__i18__net5 26.7741
rl138 n314__i18__net5 n315__i18__net5 29.8991
rl139 n320__i18__net5 n321__i18__net5 26.7741
rl140 n321__i18__net5 n322__i18__net5 29.8991
rl141 n325__i18__net5 n326__i18__net5 26.7741
rl142 n326__i18__net5 n327__i18__net5 29.8991
rl143 n328__i18__net5 n329__i18__net5 26.7741
rl144 n329__i18__net5 n330__i18__net5 29.8991
rl145 n335__i18__net5 n336__i18__net5 26.7741
rl146 n336__i18__net5 n337__i18__net5 29.8991
rl147 n338__i18__net5 n339__i18__net5 26.7741
rl148 n339__i18__net5 n340__i18__net5 29.8991
rl149 n345__i18__net5 n346__i18__net5 26.7741
rl150 n346__i18__net5 n347__i18__net5 29.8991
rl151 n348__i18__net5 n349__i18__net5 26.7741
rl152 n349__i18__net5 n350__i18__net5 29.8991
rl153 n1__ck n2__ck 202.615
rl154 n2__ck n3__ck 33.3841
rl155 n1__reset n2__reset 152.615
rl156 n2__reset n3__reset 83.3841
rl157 i14__net9 n2__i14__net9 126.36
rl158 i14__net10 n2__i14__net10 87.898
rl159 n3__i14__net10 n4__i14__net10 87.898
rl160 n3__i14__net9 n4__i14__net9 126.36
rl161 n5__i14__net9 n6__i14__net9 126.36
rl162 n5__i14__net10 n6__i14__net10 87.898
rl163 n7__i14__net10 n8__i14__net10 87.898
rl164 n7__i14__net9 n8__i14__net9 126.36
rl165 n355__i18__net5 n356__i18__net5 26.7741
rl166 n356__i18__net5 n357__i18__net5 29.8991
rl167 i14__i17__net3 n2__i14__i17__net3 126.36
rl168 n4__ck n5__ck 87.898
rl169 i14__i17__net7 n2__i14__i17__net7 87.898
rl170 i14__i17__net1 n2__i14__i17__net1 126.36
rl171 n360__i18__net5 n361__i18__net5 26.7741
rl172 n361__i18__net5 n362__i18__net5 29.8991
rl173 i14__i13__net2 n2__i14__i13__net2 11.2742
rl174 i14__i13__net2 n3__i14__i13__net2 9.7184
rl175 i14__i16__net2 n2__i14__i16__net2 9.7184
rl176 i14__i16__net2 n3__i14__i16__net2 11.2742
rl177 i14__i10__net2 n2__i14__i10__net2 11.2742
rl178 i14__i10__net2 n3__i14__i10__net2 9.7184
rl179 i14__i9__net2 n2__i14__i9__net2 9.7184
rl180 i14__i9__net2 n3__i14__i9__net2 11.2742
rl181 n365__i18__net5 n366__i18__net5 26.7741
rl182 n366__i18__net5 n367__i18__net5 29.8991
rl183 n368__i18__net5 n369__i18__net5 26.7741
rl184 n369__i18__net5 n370__i18__net5 29.8991
rl185 i14__i17__i2__net2 n2__i14__i17__i2__net2 11.2742
rl186 i14__i17__i2__net2 n3__i14__i17__i2__net2 9.7184
rl187 i14__i17__i3__net2 n2__i14__i17__i3__net2 9.7184
rl188 i14__i17__i3__net2 n3__i14__i17__i3__net2 11.2742
rl189 i14__net3 n2__i14__net3 98.1035
rl190 n3__i14__net3 n4__i14__net3 98.1035
rl191 n5__i14__net3 n6__i14__net3 98.1035
rl192 n7__i14__net3 n8__i14__net3 98.1035
rl193 n375__i18__net5 n376__i18__net5 26.7741
rl194 n376__i18__net5 n377__i18__net5 29.8991
rl195 n4__reset n5__reset 98.1035
rl196 n6__reset n7__reset 98.1035
rl197 n378__i18__net5 n379__i18__net5 26.7741
rl198 n379__i18__net5 n380__i18__net5 29.8991
rl199 i14__i13__net1 n2__i14__i13__net1 56.5719
rl200 n2__i14__i13__net1 n3__i14__i13__net1 23.6889
rl201 n3__i14__i13__net1 n4__i14__i13__net1 50.6296
rl202 n2__i14__i13__net1 n5__i14__i13__net1 56.5719
rl203 n3__i14__i13__net1 n6__i14__i13__net1 55.6157
rl204 n3__i14__i13__net1 n7__i14__i13__net1 55.6157
rl205 i14__i16__net1 n2__i14__i16__net1 56.5719
rl206 n2__i14__i16__net1 n3__i14__i16__net1 23.6889
rl207 n3__i14__i16__net1 n4__i14__i16__net1 50.6296
rl208 n2__i14__i16__net1 n5__i14__i16__net1 56.5719
rl209 n3__i14__i16__net1 n6__i14__i16__net1 55.6157
rl210 n3__i14__i16__net1 n7__i14__i16__net1 55.6157
rl211 i14__i10__net1 n2__i14__i10__net1 56.5719
rl212 n2__i14__i10__net1 n3__i14__i10__net1 23.6889
rl213 n3__i14__i10__net1 n4__i14__i10__net1 50.6296
rl214 n2__i14__i10__net1 n5__i14__i10__net1 56.5719
rl215 n3__i14__i10__net1 n6__i14__i10__net1 55.6157
rl216 n3__i14__i10__net1 n7__i14__i10__net1 55.6157
rl217 i14__i9__net1 n2__i14__i9__net1 56.5719
rl218 n2__i14__i9__net1 n3__i14__i9__net1 23.6889
rl219 n3__i14__i9__net1 n4__i14__i9__net1 50.6296
rl220 n2__i14__i9__net1 n5__i14__i9__net1 56.5719
rl221 n3__i14__i9__net1 n6__i14__i9__net1 55.6157
rl222 n3__i14__i9__net1 n7__i14__i9__net1 55.6157
rl223 n385__i18__net5 n386__i18__net5 26.7741
rl224 n386__i18__net5 n387__i18__net5 29.8991
rl225 i14__i17__i2__net1 n2__i14__i17__i2__net1 56.5719
rl226 n2__i14__i17__i2__net1 n3__i14__i17__i2__net1 23.6889
rl227 n3__i14__i17__i2__net1 n4__i14__i17__i2__net1 50.6296
rl228 n2__i14__i17__i2__net1 n5__i14__i17__i2__net1 56.5719
rl229 n3__i14__i17__i2__net1 n6__i14__i17__i2__net1 55.6157
rl230 n3__i14__i17__i2__net1 n7__i14__i17__i2__net1 55.6157
rl231 i14__i17__i3__net1 n2__i14__i17__i3__net1 56.5719
rl232 n2__i14__i17__i3__net1 n3__i14__i17__i3__net1 23.6889
rl233 n3__i14__i17__i3__net1 n4__i14__i17__i3__net1 50.6296
rl234 n2__i14__i17__i3__net1 n5__i14__i17__i3__net1 56.5719
rl235 n3__i14__i17__i3__net1 n6__i14__i17__i3__net1 55.6157
rl236 n3__i14__i17__i3__net1 n7__i14__i17__i3__net1 55.6157
rl237 n9__i14__net10 n10__i14__net10 126.36
rl238 n9__i14__net9 n10__i14__net9 87.898
rl239 n11__i14__net9 n12__i14__net9 87.898
rl240 n11__i14__net10 n12__i14__net10 126.36
rl241 n13__i14__net10 n14__i14__net10 126.36
rl242 n13__i14__net9 n14__i14__net9 87.898
rl243 n15__i14__net9 n16__i14__net9 87.898
rl244 n15__i14__net10 n16__i14__net10 126.36
rl245 n390__i18__net5 n391__i18__net5 26.7741
rl246 n391__i18__net5 n392__i18__net5 29.8991
rl247 n395__i18__net5 n396__i18__net5 26.7741
rl248 n396__i18__net5 n397__i18__net5 29.8991
rl249 n6__ck n7__ck 126.36
rl250 n3__i14__i17__net3 n4__i14__i17__net3 87.898
rl251 n3__i14__i17__net1 n4__i14__i17__net1 87.898
rl252 n3__i14__i17__net7 n4__i14__i17__net7 126.36
rl253 n398__i18__net5 n399__i18__net5 26.7741
rl254 n399__i18__net5 n400__i18__net5 29.8991
rl255 i14__i13__net4 n2__i14__i13__net4 11.2742
rl256 i14__i13__net4 n3__i14__i13__net4 9.7184
rl257 i14__i16__net4 n2__i14__i16__net4 9.7184
rl258 i14__i16__net4 n3__i14__i16__net4 11.2742
rl259 i14__i10__net4 n2__i14__i10__net4 11.2742
rl260 i14__i10__net4 n3__i14__i10__net4 9.7184
rl261 i14__i9__net4 n2__i14__i9__net4 9.7184
rl262 i14__i9__net4 n3__i14__i9__net4 11.2742
rl263 i14__net4 n2__i14__net4 74.5009
rl264 n3__i14__net4 n4__i14__net4 74.5009
rl265 n5__i14__net4 n6__i14__net4 74.5009
rl266 n7__i14__net4 n8__i14__net4 74.5009
rl267 n405__i18__net5 n406__i18__net5 26.7741
rl268 n406__i18__net5 n407__i18__net5 29.8991
rl269 i14__i17__i2__net4 n2__i14__i17__i2__net4 11.2742
rl270 i14__i17__i2__net4 n3__i14__i17__i2__net4 9.7184
rl271 i14__i17__i3__net4 n2__i14__i17__i3__net4 9.7184
rl272 i14__i17__i3__net4 n3__i14__i17__i3__net4 11.2742
rl273 n408__i18__net5 n409__i18__net5 26.7741
rl274 n409__i18__net5 n410__i18__net5 29.8991
rl275 i14__i17__net6 n2__i14__i17__net6 74.5009
rl276 n3__i14__i17__net6 n4__i14__i17__net6 74.5009
rl277 i14__i13__net5 n2__i14__i13__net5 56.5719
rl278 n2__i14__i13__net5 n3__i14__i13__net5 23.6889
rl279 n3__i14__i13__net5 n4__i14__i13__net5 50.6296
rl280 n2__i14__i13__net5 n5__i14__i13__net5 56.5719
rl281 n3__i14__i13__net5 n6__i14__i13__net5 55.6157
rl282 n3__i14__i13__net5 n7__i14__i13__net5 55.6157
rl283 i14__i16__net5 n2__i14__i16__net5 56.5719
rl284 n2__i14__i16__net5 n3__i14__i16__net5 23.6889
rl285 n3__i14__i16__net5 n4__i14__i16__net5 50.6296
rl286 n2__i14__i16__net5 n5__i14__i16__net5 56.5719
rl287 n3__i14__i16__net5 n6__i14__i16__net5 55.6157
rl288 n3__i14__i16__net5 n7__i14__i16__net5 55.6157
rl289 i14__i10__net5 n2__i14__i10__net5 56.5719
rl290 n2__i14__i10__net5 n3__i14__i10__net5 23.6889
rl291 n3__i14__i10__net5 n4__i14__i10__net5 50.6296
rl292 n2__i14__i10__net5 n5__i14__i10__net5 56.5719
rl293 n3__i14__i10__net5 n6__i14__i10__net5 55.6157
rl294 n3__i14__i10__net5 n7__i14__i10__net5 55.6157
rl295 i14__i9__net5 n2__i14__i9__net5 56.5719
rl296 n2__i14__i9__net5 n3__i14__i9__net5 23.6889
rl297 n3__i14__i9__net5 n4__i14__i9__net5 50.6296
rl298 n2__i14__i9__net5 n5__i14__i9__net5 56.5719
rl299 n3__i14__i9__net5 n6__i14__i9__net5 55.6157
rl300 n3__i14__i9__net5 n7__i14__i9__net5 55.6157
rl301 n413__i18__net5 n414__i18__net5 26.7741
rl302 n414__i18__net5 n415__i18__net5 29.8991
rl303 n4__i14__i13__net4 n5__i14__i13__net4 49.0903
rl304 n5__i14__i13__net4 n6__i14__i13__net4 49.0903
rl305 n4__i14__i16__net4 n5__i14__i16__net4 49.0903
rl306 n5__i14__i16__net4 n6__i14__i16__net4 49.0903
rl307 n4__i14__i10__net4 n5__i14__i10__net4 49.0903
rl308 n5__i14__i10__net4 n6__i14__i10__net4 49.0903
rl309 n4__i14__i9__net4 n5__i14__i9__net4 49.0903
rl310 n5__i14__i9__net4 n6__i14__i9__net4 49.0903
rl311 i14__i17__i2__net5 n2__i14__i17__i2__net5 56.5719
rl312 n2__i14__i17__i2__net5 n3__i14__i17__i2__net5 23.6889
rl313 n3__i14__i17__i2__net5 n4__i14__i17__i2__net5 50.6296
rl314 n2__i14__i17__i2__net5 n5__i14__i17__i2__net5 56.5719
rl315 n3__i14__i17__i2__net5 n6__i14__i17__i2__net5 55.6157
rl316 n3__i14__i17__i2__net5 n7__i14__i17__i2__net5 55.6157
rl317 i14__i17__i3__net5 n2__i14__i17__i3__net5 56.5719
rl318 n2__i14__i17__i3__net5 n3__i14__i17__i3__net5 23.6889
rl319 n3__i14__i17__i3__net5 n4__i14__i17__i3__net5 50.6296
rl320 n2__i14__i17__i3__net5 n5__i14__i17__i3__net5 56.5719
rl321 n3__i14__i17__i3__net5 n6__i14__i17__i3__net5 55.6157
rl322 n3__i14__i17__i3__net5 n7__i14__i17__i3__net5 55.6157
rl323 n419__i18__net5 n420__i18__net5 26.7741
rl324 n420__i18__net5 n421__i18__net5 29.8991
rl325 n423__i18__net5 n424__i18__net5 26.7741
rl326 n424__i18__net5 n425__i18__net5 29.8991
rl327 i14__y_out_b_3 n2__i14__y_out_b_3 56.5719
rl328 n2__i14__y_out_b_3 n3__i14__y_out_b_3 50.013
rl329 n2__i14__y_out_b_3 n4__i14__y_out_b_3 56.5719
rl330 i14__y_out_b_0 n2__i14__y_out_b_0 56.5719
rl331 n2__i14__y_out_b_0 n3__i14__y_out_b_0 50.013
rl332 n2__i14__y_out_b_0 n4__i14__y_out_b_0 56.5719
rl333 i14__x_out_b_2 n2__i14__x_out_b_2 56.5719
rl334 n2__i14__x_out_b_2 n3__i14__x_out_b_2 50.013
rl335 n2__i14__x_out_b_2 n4__i14__x_out_b_2 56.5719
rl336 i14__x_out_b_3 n2__i14__x_out_b_3 56.5719
rl337 n2__i14__x_out_b_3 n3__i14__x_out_b_3 50.013
rl338 n2__i14__x_out_b_3 n4__i14__x_out_b_3 56.5719
rl339 n4__i14__i17__i2__net4 n5__i14__i17__i2__net4 49.0903
rl340 n5__i14__i17__i2__net4 n6__i14__i17__i2__net4 49.0903
rl341 n4__i14__i17__i3__net4 n5__i14__i17__i3__net4 49.0903
rl342 n5__i14__i17__i3__net4 n6__i14__i17__i3__net4 49.0903
rl343 n428__i18__net5 n429__i18__net5 26.7741
rl344 n429__i18__net5 n430__i18__net5 29.8991
rl345 n14__i14__i17__net1 n15__i14__i17__net1 56.5719
rl346 n15__i14__i17__net1 n16__i14__i17__net1 50.013
rl347 n15__i14__i17__net1 n17__i14__i17__net1 56.5719
rl348 n6__i14__i17__net8 n7__i14__i17__net8 56.5719
rl349 n7__i14__i17__net8 n8__i14__i17__net8 50.013
rl350 n7__i14__i17__net8 n9__i14__i17__net8 56.5719
rl351 n33__i14__net9 n34__i14__net9 126.36
rl352 n29__i14__net10 n30__i14__net10 87.898
rl353 n31__i14__net10 n32__i14__net10 87.898
rl354 n35__i14__net9 n36__i14__net9 126.36
rl355 n37__i14__net9 n38__i14__net9 126.36
rl356 n33__i14__net10 n34__i14__net10 87.898
rl357 n35__i14__net10 n36__i14__net10 87.898
rl358 n39__i14__net9 n40__i14__net9 126.36
rl359 n435__i18__net5 n436__i18__net5 26.7741
rl360 n436__i18__net5 n437__i18__net5 29.8991
rl361 i14__i17__net10 n2__i14__i17__net10 56.5719
rl362 n2__i14__i17__net10 n3__i14__i17__net10 48.1183
rl363 n2__i14__i17__net10 n4__i14__i17__net10 56.5719
rl364 n10__i14__i17__net8 n11__i14__i17__net8 69.2328
rl365 n440__i18__net5 n441__i18__net5 26.7741
rl366 n441__i18__net5 n442__i18__net5 29.8991
rl367 i14__i17__net11 n2__i14__i17__net11 101.925
rl368 n2__i14__i17__net11 n3__i14__i17__net11 201.489
rl369 n12__i14__i17__net8 n13__i14__i17__net8 73.079
rl370 n443__i18__net5 n444__i18__net5 26.7741
rl371 n444__i18__net5 n445__i18__net5 29.8991
rl372 i14__i17__net9 n2__i14__i17__net9 56.5719
rl373 n2__i14__i17__net9 n3__i14__i17__net9 48.1183
rl374 n2__i14__i17__net9 n4__i14__i17__net9 56.5719
rl375 i14__i11__net2 n2__i14__i11__net2 11.2742
rl376 i14__i11__net2 n3__i14__i11__net2 9.7184
rl377 i14__i14__net2 n2__i14__i14__net2 9.7184
rl378 i14__i14__net2 n3__i14__i14__net2 11.2742
rl379 i14__i15__net2 n2__i14__i15__net2 11.2742
rl380 i14__i15__net2 n3__i14__i15__net2 9.7184
rl381 i14__i12__net2 n2__i14__i12__net2 9.7184
rl382 i14__i12__net2 n3__i14__i12__net2 11.2742
rl383 n5__i14__i17__net9 n6__i14__i17__net9 64.1533
rl384 n6__i14__i17__net9 n7__i14__i17__net9 33.3841
rl385 n450__i18__net5 n451__i18__net5 26.7741
rl386 n451__i18__net5 n452__i18__net5 29.8991
rl387 n453__i18__net5 n454__i18__net5 26.7741
rl388 n454__i18__net5 n455__i18__net5 29.8991
rl389 n29__i14__net3 n30__i14__net3 98.1035
rl390 n31__i14__net3 n32__i14__net3 98.1035
rl391 n33__i14__net3 n34__i14__net3 98.1035
rl392 n35__i14__net3 n36__i14__net3 98.1035
rl393 n5__i14__i17__net10 n6__i14__i17__net10 33.3841
rl394 n6__i14__i17__net10 n7__i14__i17__net10 64.1533
rl395 n458__i18__net5 n459__i18__net5 26.7741
rl396 n459__i18__net5 n460__i18__net5 29.8991
rl397 n4__i14__i17__net11 n5__i14__i17__net11 73.079
rl398 i14__i11__net1 n2__i14__i11__net1 56.5719
rl399 n2__i14__i11__net1 n3__i14__i11__net1 23.6889
rl400 n3__i14__i11__net1 n4__i14__i11__net1 50.6296
rl401 n2__i14__i11__net1 n5__i14__i11__net1 56.5719
rl402 n3__i14__i11__net1 n6__i14__i11__net1 55.6157
rl403 n3__i14__i11__net1 n7__i14__i11__net1 55.6157
rl404 i14__i14__net1 n2__i14__i14__net1 56.5719
rl405 n2__i14__i14__net1 n3__i14__i14__net1 23.6889
rl406 n3__i14__i14__net1 n4__i14__i14__net1 50.6296
rl407 n2__i14__i14__net1 n5__i14__i14__net1 56.5719
rl408 n3__i14__i14__net1 n6__i14__i14__net1 55.6157
rl409 n3__i14__i14__net1 n7__i14__i14__net1 55.6157
rl410 i14__i15__net1 n2__i14__i15__net1 56.5719
rl411 n2__i14__i15__net1 n3__i14__i15__net1 23.6889
rl412 n3__i14__i15__net1 n4__i14__i15__net1 50.6296
rl413 n2__i14__i15__net1 n5__i14__i15__net1 56.5719
rl414 n3__i14__i15__net1 n6__i14__i15__net1 55.6157
rl415 n3__i14__i15__net1 n7__i14__i15__net1 55.6157
rl416 i14__i12__net1 n2__i14__i12__net1 56.5719
rl417 n2__i14__i12__net1 n3__i14__i12__net1 23.6889
rl418 n3__i14__i12__net1 n4__i14__i12__net1 50.6296
rl419 n2__i14__i12__net1 n5__i14__i12__net1 56.5719
rl420 n3__i14__i12__net1 n6__i14__i12__net1 55.6157
rl421 n3__i14__i12__net1 n7__i14__i12__net1 55.6157
rl422 n463__i18__net5 n464__i18__net5 26.7741
rl423 n464__i18__net5 n465__i18__net5 29.8991
rl424 n14__i14__i17__net8 n15__i14__i17__net8 201.489
rl425 n15__i14__i17__net8 n16__i14__i17__net8 69.2328
rl426 n6__i14__i17__net11 n7__i14__i17__net11 101.925
rl427 n26__reset n27__reset 56.5719
rl428 n27__reset n28__reset 23.6889
rl429 n28__reset n29__reset 10.1559
rl430 n29__reset n30__reset 8.8401
rl431 n30__reset n31__reset 26.2002
rl432 n31__reset n32__reset 9.498
rl433 n32__reset n33__reset 9.498
rl434 n33__reset n34__reset 23.6922
rl435 n34__reset n35__reset 56.5719
rl436 n27__reset n36__reset 56.5719
rl437 n28__reset n37__reset 55.6157
rl438 n28__reset n38__reset 55.6157
rl439 n30__reset n39__reset 55.6157
rl440 n30__reset n40__reset 55.6157
rl441 n31__reset n41__reset 55.6157
rl442 n31__reset n42__reset 55.6157
rl443 n33__reset n43__reset 55.6157
rl444 n33__reset n44__reset 55.6157
rl445 n34__reset n45__reset 56.5719
rl446 n470__i18__net5 n471__i18__net5 24.7396
rl447 n471__i18__net5 n472__i18__net5 23.2442
rl448 n57__i14__net10 n58__i14__net10 126.36
rl449 n49__i14__net9 n50__i14__net9 87.898
rl450 n51__i14__net9 n52__i14__net9 87.898
rl451 n59__i14__net10 n60__i14__net10 126.36
rl452 n61__i14__net10 n62__i14__net10 126.36
rl453 n53__i14__net9 n54__i14__net9 87.898
rl454 n55__i14__net9 n56__i14__net9 87.898
rl455 n63__i14__net10 n64__i14__net10 126.36
rl456 i14__net7 n2__i14__net7 56.5719
rl457 n2__i14__net7 n3__i14__net7 48.1183
rl458 n2__i14__net7 n4__i14__net7 56.5719
rl459 i14__i11__net4 n2__i14__i11__net4 11.2742
rl460 i14__i11__net4 n3__i14__i11__net4 9.7184
rl461 i14__i14__net4 n2__i14__i14__net4 9.7184
rl462 i14__i14__net4 n3__i14__i14__net4 11.2742
rl463 i14__i15__net4 n2__i14__i15__net4 11.2742
rl464 i14__i15__net4 n3__i14__i15__net4 9.7184
rl465 i14__i12__net4 n2__i14__i12__net4 9.7184
rl466 i14__i12__net4 n3__i14__i12__net4 11.2742
rl467 n21__i14__net4 n22__i14__net4 74.5009
rl468 n23__i14__net4 n24__i14__net4 74.5009
rl469 n25__i14__net4 n26__i14__net4 74.5009
rl470 n27__i14__net4 n28__i14__net4 74.5009
rl471 i14__net11 n2__i14__net11 56.5719
rl472 n2__i14__net11 n3__i14__net11 48.1183
rl473 n2__i14__net11 n4__i14__net11 56.5719
rl474 n29__i14__net4 n30__i14__net4 56.5719
rl475 n30__i14__net4 n31__i14__net4 23.6889
rl476 n31__i14__net4 n32__i14__net4 9.498
rl477 n32__i14__net4 n33__i14__net4 9.498
rl478 n33__i14__net4 n34__i14__net4 26.2002
rl479 n34__i14__net4 n35__i14__net4 9.498
rl480 n35__i14__net4 n36__i14__net4 9.498
rl481 n36__i14__net4 n37__i14__net4 23.6922
rl482 n37__i14__net4 n38__i14__net4 56.5719
rl483 n30__i14__net4 n39__i14__net4 56.5719
rl484 n31__i14__net4 n40__i14__net4 55.6157
rl485 n31__i14__net4 n41__i14__net4 55.6157
rl486 n33__i14__net4 n42__i14__net4 55.6157
rl487 n33__i14__net4 n43__i14__net4 55.6157
rl488 n34__i14__net4 n44__i14__net4 55.6157
rl489 n34__i14__net4 n45__i14__net4 55.6157
rl490 n36__i14__net4 n46__i14__net4 55.6157
rl491 n36__i14__net4 n47__i14__net4 55.6157
rl492 n37__i14__net4 n48__i14__net4 56.5719
rl493 i14__i11__net5 n2__i14__i11__net5 56.5719
rl494 n2__i14__i11__net5 n3__i14__i11__net5 23.6889
rl495 n3__i14__i11__net5 n4__i14__i11__net5 50.6296
rl496 n2__i14__i11__net5 n5__i14__i11__net5 56.5719
rl497 n3__i14__i11__net5 n6__i14__i11__net5 55.6157
rl498 n3__i14__i11__net5 n7__i14__i11__net5 55.6157
rl499 i14__i14__net5 n2__i14__i14__net5 56.5719
rl500 n2__i14__i14__net5 n3__i14__i14__net5 23.6889
rl501 n3__i14__i14__net5 n4__i14__i14__net5 50.6296
rl502 n2__i14__i14__net5 n5__i14__i14__net5 56.5719
rl503 n3__i14__i14__net5 n6__i14__i14__net5 55.6157
rl504 n3__i14__i14__net5 n7__i14__i14__net5 55.6157
rl505 i14__i15__net5 n2__i14__i15__net5 56.5719
rl506 n2__i14__i15__net5 n3__i14__i15__net5 23.6889
rl507 n3__i14__i15__net5 n4__i14__i15__net5 50.6296
rl508 n2__i14__i15__net5 n5__i14__i15__net5 56.5719
rl509 n3__i14__i15__net5 n6__i14__i15__net5 55.6157
rl510 n3__i14__i15__net5 n7__i14__i15__net5 55.6157
rl511 i14__i12__net5 n2__i14__i12__net5 56.5719
rl512 n2__i14__i12__net5 n3__i14__i12__net5 23.6889
rl513 n3__i14__i12__net5 n4__i14__i12__net5 50.6296
rl514 n2__i14__i12__net5 n5__i14__i12__net5 56.5719
rl515 n3__i14__i12__net5 n6__i14__i12__net5 55.6157
rl516 n3__i14__i12__net5 n7__i14__i12__net5 55.6157
rl517 i18__net4 n2__i18__net4 26.7741
rl518 n2__i18__net4 n3__i18__net4 29.8991
rl519 n4__i14__i11__net4 n5__i14__i11__net4 49.0903
rl520 n5__i14__i11__net4 n6__i14__i11__net4 49.0903
rl521 n4__i14__i14__net4 n5__i14__i14__net4 49.0903
rl522 n5__i14__i14__net4 n6__i14__i14__net4 49.0903
rl523 n4__i14__i15__net4 n5__i14__i15__net4 49.0903
rl524 n5__i14__i15__net4 n6__i14__i15__net4 49.0903
rl525 n4__i14__i12__net4 n5__i14__i12__net4 49.0903
rl526 n5__i14__i12__net4 n6__i14__i12__net4 49.0903
rl527 n4__i18__net4 n5__i18__net4 26.7741
rl528 n5__i18__net4 n6__i18__net4 29.8991
rl529 n7__i18__net4 n8__i18__net4 26.7741
rl530 n8__i18__net4 n9__i18__net4 29.8991
rl531 n5__i14__net7 n6__i14__net7 56.5719
rl532 n6__i14__net7 n7__i14__net7 23.6889
rl533 n7__i14__net7 n8__i14__net7 9.498
rl534 n8__i14__net7 n9__i14__net7 9.498
rl535 n9__i14__net7 n10__i14__net7 26.2002
rl536 n10__i14__net7 n11__i14__net7 9.498
rl537 n11__i14__net7 n12__i14__net7 9.498
rl538 n12__i14__net7 n13__i14__net7 23.6922
rl539 n13__i14__net7 n14__i14__net7 56.5719
rl540 n6__i14__net7 n15__i14__net7 56.5719
rl541 n7__i14__net7 n16__i14__net7 55.6157
rl542 n7__i14__net7 n17__i14__net7 55.6157
rl543 n9__i14__net7 n18__i14__net7 55.6157
rl544 n9__i14__net7 n19__i14__net7 55.6157
rl545 n10__i14__net7 n20__i14__net7 55.6157
rl546 n10__i14__net7 n21__i14__net7 55.6157
rl547 n12__i14__net7 n22__i14__net7 55.6157
rl548 n12__i14__net7 n23__i14__net7 55.6157
rl549 n13__i14__net7 n24__i14__net7 56.5719
rl550 n5__i14__net11 n6__i14__net11 56.5719
rl551 n6__i14__net11 n7__i14__net11 23.6889
rl552 n7__i14__net11 n8__i14__net11 9.498
rl553 n8__i14__net11 n9__i14__net11 9.498
rl554 n9__i14__net11 n10__i14__net11 26.2002
rl555 n10__i14__net11 n11__i14__net11 9.498
rl556 n11__i14__net11 n12__i14__net11 9.498
rl557 n12__i14__net11 n13__i14__net11 23.6922
rl558 n13__i14__net11 n14__i14__net11 56.5719
rl559 n6__i14__net11 n15__i14__net11 56.5719
rl560 n7__i14__net11 n16__i14__net11 55.6157
rl561 n7__i14__net11 n17__i14__net11 55.6157
rl562 n9__i14__net11 n18__i14__net11 55.6157
rl563 n9__i14__net11 n19__i14__net11 55.6157
rl564 n10__i14__net11 n20__i14__net11 55.6157
rl565 n10__i14__net11 n21__i14__net11 55.6157
rl566 n12__i14__net11 n22__i14__net11 55.6157
rl567 n12__i14__net11 n23__i14__net11 55.6157
rl568 n13__i14__net11 n24__i14__net11 56.5719
rl569 i14__x_out_b_1 n2__i14__x_out_b_1 56.5719
rl570 n2__i14__x_out_b_1 n3__i14__x_out_b_1 50.013
rl571 n2__i14__x_out_b_1 n4__i14__x_out_b_1 56.5719
rl572 i14__y_out_b_2 n2__i14__y_out_b_2 56.5719
rl573 n2__i14__y_out_b_2 n3__i14__y_out_b_2 50.013
rl574 n2__i14__y_out_b_2 n4__i14__y_out_b_2 56.5719
rl575 i14__y_out_b_1 n2__i14__y_out_b_1 56.5719
rl576 n2__i14__y_out_b_1 n3__i14__y_out_b_1 50.013
rl577 n2__i14__y_out_b_1 n4__i14__y_out_b_1 56.5719
rl578 i14__x_out_b_0 n2__i14__x_out_b_0 56.5719
rl579 n2__i14__x_out_b_0 n3__i14__x_out_b_0 50.013
rl580 n2__i14__x_out_b_0 n4__i14__x_out_b_0 56.5719
rl581 n10__i18__net4 n11__i18__net4 26.7741
rl582 n11__i18__net4 n12__i18__net4 29.8991
rl583 n13__i18__net4 n14__i18__net4 26.7741
rl584 n14__i18__net4 n15__i18__net4 29.8991
rl585 n6__x_out_2 n7__x_out_2 56.5719
rl586 n7__x_out_2 n8__x_out_2 48.1183
rl587 n7__x_out_2 n9__x_out_2 56.5719
rl588 y_out_0 n2__y_out_0 56.5719
rl589 n2__y_out_0 n3__y_out_0 48.1183
rl590 n2__y_out_0 n4__y_out_0 56.5719
rl591 ck_buff n2__ck_buff 87.898
rl592 ck_b n2__ck_b 126.36
rl593 n16__i18__net4 n17__i18__net4 26.7741
rl594 n17__i18__net4 n18__i18__net4 29.8991
rl595 n10__x_out_2 n11__x_out_2 87.2876
rl596 n5__y_out_0 n6__y_out_0 87.2876
rl597 i13__i14__net2 n2__i13__i14__net2 82.6365
rl598 i13__i12__net2 n2__i13__i12__net2 82.6365
rl599 net11 n2__net11 45
rl600 n2__net11 n3__net11 26.2002
rl601 n3__net11 n4__net11 20.3369
rl602 n2__net11 n5__net11 55.6157
rl603 n2__net11 n6__net11 55.6157
rl604 n3__net11 n7__net11 55.6157
rl605 n3__net11 n8__net11 55.6157
rl606 n4__net11 n9__net11 47.7829
rl607 n4__net11 n10__net11 47.7829
rl608 n19__i18__net4 n20__i18__net4 26.7741
rl609 n20__i18__net4 n21__i18__net4 29.8991
rl610 y_out_2 n2__y_out_2 56.5719
rl611 n2__y_out_2 n3__y_out_2 48.1183
rl612 n2__y_out_2 n4__y_out_2 56.5719
rl613 n6__x_out_0 n7__x_out_0 56.5719
rl614 n7__x_out_0 n8__x_out_0 48.1183
rl615 n7__x_out_0 n9__x_out_0 56.5719
rl616 n22__i18__net4 n23__i18__net4 26.7741
rl617 n23__i18__net4 n24__i18__net4 29.8991
rl618 i9__i4__net2 n2__i9__i4__net2 9.7184
rl619 i9__i4__net2 n3__i9__i4__net2 11.2742
rl620 n25__i18__net4 n26__i18__net4 26.7741
rl621 n26__i18__net4 n27__i18__net4 29.8991
rl622 net9 n2__net9 45
rl623 n2__net9 n3__net9 26.2002
rl624 n3__net9 n4__net9 23.6922
rl625 n4__net9 n5__net9 56.5719
rl626 n2__net9 n6__net9 55.6157
rl627 n2__net9 n7__net9 55.6157
rl628 n3__net9 n8__net9 55.6157
rl629 n3__net9 n9__net9 55.6157
rl630 n4__net9 n10__net9 56.5719
rl631 n28__i18__net4 n29__i18__net4 26.7741
rl632 n29__i18__net4 n30__i18__net4 29.8991
rl633 reset_buff n2__reset_buff 98.1035
rl634 n31__i18__net4 n32__i18__net4 26.7741
rl635 n32__i18__net4 n33__i18__net4 29.8991
rl636 n6__x_out_3 n7__x_out_3 56.5719
rl637 n7__x_out_3 n8__x_out_3 48.1183
rl638 n7__x_out_3 n9__x_out_3 56.5719
rl639 n6__x_out_1 n7__x_out_1 56.5719
rl640 n7__x_out_1 n8__x_out_1 48.1183
rl641 n7__x_out_1 n9__x_out_1 56.5719
rl642 n22__ck n23__ck 45
rl643 n23__ck n24__ck 56.5719
rl644 n23__ck n25__ck 56.5719
rl645 i9__i4__net1 n2__i9__i4__net1 56.5719
rl646 n2__i9__i4__net1 n3__i9__i4__net1 23.6889
rl647 n3__i9__i4__net1 n4__i9__i4__net1 50.6296
rl648 n2__i9__i4__net1 n5__i9__i4__net1 56.5719
rl649 n3__i9__i4__net1 n6__i9__i4__net1 55.6157
rl650 n3__i9__i4__net1 n7__i9__i4__net1 55.6157
rl651 n34__i18__net4 n35__i18__net4 26.7741
rl652 n35__i18__net4 n36__i18__net4 29.8991
rl653 n10__x_out_3 n11__x_out_3 87.2876
rl654 n10__x_out_1 n11__x_out_1 87.2876
rl655 i13__i15__net2 n2__i13__i15__net2 82.6365
rl656 i13__i13__net2 n2__i13__i13__net2 82.6365
rl657 n37__i18__net4 n38__i18__net4 26.7741
rl658 n38__i18__net4 n39__i18__net4 29.8991
rl659 n3__ck_b n4__ck_b 87.898
rl660 n3__ck_buff n4__ck_buff 126.36
rl661 net12 n2__net12 45
rl662 n2__net12 n3__net12 26.2002
rl663 n3__net12 n4__net12 20.3369
rl664 n2__net12 n5__net12 55.6157
rl665 n2__net12 n6__net12 55.6157
rl666 n3__net12 n7__net12 55.6157
rl667 n3__net12 n8__net12 55.6157
rl668 n4__net12 n9__net12 47.7829
rl669 n4__net12 n10__net12 47.7829
rl670 n40__i18__net4 n41__i18__net4 26.7741
rl671 n41__i18__net4 n42__i18__net4 29.8991
rl672 y_out_3 n2__y_out_3 56.5719
rl673 n2__y_out_3 n3__y_out_3 48.1183
rl674 n2__y_out_3 n4__y_out_3 56.5719
rl675 y_out_1 n2__y_out_1 56.5719
rl676 n2__y_out_1 n3__y_out_1 48.1183
rl677 n2__y_out_1 n4__y_out_1 56.5719
rl678 n45__i18__net4 n46__i18__net4 26.7741
rl679 n46__i18__net4 n47__i18__net4 29.8991
rl680 i9__i4__net4 n2__i9__i4__net4 9.7184
rl681 i9__i4__net4 n3__i9__i4__net4 11.2742
rl682 n48__i18__net4 n49__i18__net4 26.7741
rl683 n49__i18__net4 n50__i18__net4 29.8991
rl684 reset_b n2__reset_b 74.5009
rl685 net10 n2__net10 45
rl686 n2__net10 n3__net10 26.2002
rl687 n3__net10 n4__net10 23.6922
rl688 n4__net10 n5__net10 56.5719
rl689 n2__net10 n6__net10 55.6157
rl690 n2__net10 n7__net10 55.6157
rl691 n3__net10 n8__net10 55.6157
rl692 n3__net10 n9__net10 55.6157
rl693 n4__net10 n10__net10 56.5719
rl694 n53__i18__net4 n54__i18__net4 26.7741
rl695 n54__i18__net4 n55__i18__net4 29.8991
rl696 i13__a3 n2__i13__a3 137.341
rl697 n2__i13__a3 n3__i13__a3 48.1183
rl698 n2__i13__a3 n4__i13__a3 68.1104
rl699 i13__a1 n2__i13__a1 68.1104
rl700 n2__i13__a1 n3__i13__a1 48.1183
rl701 n2__i13__a1 n4__i13__a1 137.341
rl702 n26__ck n27__ck 56.5719
rl703 n27__ck n28__ck 45
rl704 n27__ck n29__ck 56.5719
rl705 i13__a2 n2__i13__a2 60.4181
rl706 n2__i13__a2 n3__i13__a2 48.1183
rl707 n2__i13__a2 n4__i13__a2 145.033
rl708 i13__a0 n2__i13__a0 145.033
rl709 n2__i13__a0 n3__i13__a0 48.1183
rl710 n2__i13__a0 n4__i13__a0 60.4181
rl711 n59__i18__net4 n60__i18__net4 26.7741
rl712 n60__i18__net4 n61__i18__net4 29.8991
rl713 n51__reset n52__reset 45
rl714 n52__reset n53__reset 56.5719
rl715 n52__reset n54__reset 56.5719
rl716 i9__i4__net5 n2__i9__i4__net5 56.5719
rl717 n2__i9__i4__net5 n3__i9__i4__net5 23.6889
rl718 n3__i9__i4__net5 n4__i9__i4__net5 50.6296
rl719 n2__i9__i4__net5 n5__i9__i4__net5 56.5719
rl720 n3__i9__i4__net5 n6__i9__i4__net5 55.6157
rl721 n3__i9__i4__net5 n7__i9__i4__net5 55.6157
rl722 n63__i18__net4 n64__i18__net4 26.7741
rl723 n64__i18__net4 n65__i18__net4 29.8991
rl724 i13__i17__net1 n2__i13__i17__net1 56.5719
rl725 n2__i13__i17__net1 n3__i13__i17__net1 48.1183
rl726 n2__i13__i17__net1 n4__i13__i17__net1 56.5719
rl727 i13__i16__net1 n2__i13__i16__net1 56.5719
rl728 n2__i13__i16__net1 n3__i13__i16__net1 48.1183
rl729 n2__i13__i16__net1 n4__i13__i16__net1 56.5719
rl730 n4__i9__i4__net4 n5__i9__i4__net4 49.0903
rl731 n5__i9__i4__net4 n6__i9__i4__net4 49.0903
rl732 n55__reset n56__reset 56.5719
rl733 n56__reset n57__reset 45
rl734 n56__reset n58__reset 56.5719
rl735 n68__i18__net4 n69__i18__net4 26.7741
rl736 n69__i18__net4 n70__i18__net4 29.8991
rl737 net13 n2__net13 48.3127
rl738 n2__net13 n3__net13 47.7829
rl739 n2__net13 n4__net13 20.3369
rl740 n4__net13 n5__net13 55.6157
rl741 n4__net13 n6__net13 26.2002
rl742 n6__net13 n7__net13 55.6157
rl743 n4__net13 n8__net13 55.6157
rl744 n6__net13 n9__net13 45
rl745 n6__net13 n10__net13 55.6157
rl746 i9__net2 n2__i9__net2 56.5719
rl747 n2__i9__net2 n3__i9__net2 50.013
rl748 n2__i9__net2 n4__i9__net2 56.5719
rl749 n5__i13__a2 n6__i13__a2 56.5719
rl750 n6__i13__a2 n7__i13__a2 48.1183
rl751 n6__i13__a2 n8__i13__a2 56.5719
rl752 n5__i13__a0 n6__i13__a0 56.5719
rl753 n6__i13__a0 n7__i13__a0 48.1183
rl754 n6__i13__a0 n8__i13__a0 56.5719
rl755 n73__i18__net4 n74__i18__net4 26.7741
rl756 n74__i18__net4 n75__i18__net4 29.8991
rl757 n80__i18__net4 n81__i18__net4 26.7741
rl758 n81__i18__net4 n82__i18__net4 29.8991
rl759 n13__i13__a2 n14__i13__a2 87.2876
rl760 n13__i13__a0 n14__i13__a0 87.2876
rl761 i13__i17__i4__net2 n2__i13__i17__i4__net2 82.6365
rl762 i13__i16__i4__net2 n2__i13__i16__i4__net2 82.6365
rl763 net14 n2__net14 48.3127
rl764 n2__net14 n3__net14 47.7829
rl765 n2__net14 n4__net14 20.3369
rl766 n4__net14 n5__net14 55.6157
rl767 n4__net14 n6__net14 26.2002
rl768 n6__net14 n7__net14 55.6157
rl769 n4__net14 n8__net14 55.6157
rl770 n6__net14 n9__net14 45
rl771 n6__net14 n10__net14 55.6157
rl772 n83__i18__net4 n84__i18__net4 26.7741
rl773 n84__i18__net4 n85__i18__net4 29.8991
rl774 i9__net1 n2__i9__net1 57.4064
rl775 n2__i9__net1 n3__i9__net1 18.4261
rl776 n2__i9__net1 n4__i9__net1 57.4064
rl777 n3__i9__net1 n5__i9__net1 49.4506
rl778 n3__i9__net1 n6__i9__net1 49.4506
rl779 n5__i13__a3 n6__i13__a3 56.5719
rl780 n6__i13__a3 n7__i13__a3 48.1183
rl781 n6__i13__a3 n8__i13__a3 56.5719
rl782 n5__i13__a1 n6__i13__a1 56.5719
rl783 n6__i13__a1 n7__i13__a1 48.1183
rl784 n6__i13__a1 n8__i13__a1 56.5719
rl785 n88__i18__net4 n89__i18__net4 26.7741
rl786 n89__i18__net4 n90__i18__net4 29.8991
rl787 n10__ck4 n11__ck4 57.4064
rl788 n11__ck4 n12__ck4 18.4261
rl789 n11__ck4 n13__ck4 57.4064
rl790 n12__ck4 n14__ck4 49.4506
rl791 n12__ck4 n15__ck4 49.4506
rl792 n95__i18__net4 n96__i18__net4 26.7741
rl793 n96__i18__net4 n97__i18__net4 29.8991
rl794 n100__i18__net4 n101__i18__net4 26.7741
rl795 n101__i18__net4 n102__i18__net4 29.8991
rl796 shift n2__shift 147.791
rl797 n2__shift n3__shift 47.7666
rl798 n2__shift n4__shift 38.1757
rl799 n5__shift n6__shift 38.1757
rl800 n6__shift n7__shift 47.7666
rl801 n6__shift n8__shift 147.791
rl802 n9__shift n10__shift 147.791
rl803 n10__shift n11__shift 47.7666
rl804 n10__shift n12__shift 38.1757
rl805 i13__net11 n2__i13__net11 137.341
rl806 n2__i13__net11 n3__i13__net11 48.1183
rl807 n2__i13__net11 n4__i13__net11 68.1104
rl808 i13__net12 n2__i13__net12 68.1104
rl809 n2__i13__net12 n3__i13__net12 48.1183
rl810 n2__i13__net12 n4__i13__net12 137.341
rl811 n103__i18__net4 n104__i18__net4 26.7741
rl812 n104__i18__net4 n105__i18__net4 29.8991
rl813 i2__net79 n2__i2__net79 78.658
rl814 n13__shift n14__shift 80.9926
rl815 n15__shift n16__shift 80.9926
rl816 i1__net79 n2__i1__net79 78.658
rl817 i0__net79 n2__i0__net79 78.658
rl818 n17__shift n18__shift 80.9926
rl819 i13__net1 n2__i13__net1 60.4181
rl820 n2__i13__net1 n3__i13__net1 48.1183
rl821 n2__i13__net1 n4__i13__net1 145.033
rl822 i13__net2 n2__i13__net2 145.033
rl823 n2__i13__net2 n3__i13__net2 48.1183
rl824 n2__i13__net2 n4__i13__net2 60.4181
rl825 n110__i18__net4 n111__i18__net4 26.7741
rl826 n111__i18__net4 n112__i18__net4 29.8991
rl827 n3__i2__net79 n4__i2__net79 75.2349
rl828 n3__i1__net79 n4__i1__net79 75.2349
rl829 n3__i0__net79 n4__i0__net79 75.2349
rl830 n19__shift n20__shift 85.9749
rl831 n21__shift n22__shift 85.9749
rl832 n23__shift n24__shift 85.9749
rl833 i13__i19__net1 n2__i13__i19__net1 56.5719
rl834 n2__i13__i19__net1 n3__i13__i19__net1 48.1183
rl835 n2__i13__i19__net1 n4__i13__i19__net1 56.5719
rl836 i13__i18__net1 n2__i13__i18__net1 56.5719
rl837 n2__i13__i18__net1 n3__i13__i18__net1 48.1183
rl838 n2__i13__i18__net1 n4__i13__i18__net1 56.5719
rl839 n113__i18__net4 n114__i18__net4 26.7741
rl840 n114__i18__net4 n115__i18__net4 29.8991
rl841 n120__i18__net4 n121__i18__net4 24.7396
rl842 n121__i18__net4 n122__i18__net4 23.2442
rl843 n5__i13__net1 n6__i13__net1 56.5719
rl844 n6__i13__net1 n7__i13__net1 48.1183
rl845 n6__i13__net1 n8__i13__net1 56.5719
rl846 n5__i13__net2 n6__i13__net2 56.5719
rl847 n6__i13__net2 n7__i13__net2 48.1183
rl848 n6__i13__net2 n8__i13__net2 56.5719
rl849 i2__net1 n2__i2__net1 56.5719
rl850 n2__i2__net1 n3__i2__net1 48.1183
rl851 n2__i2__net1 n4__i2__net1 56.5719
rl852 i1__net1 n2__i1__net1 56.5719
rl853 n2__i1__net1 n3__i1__net1 48.1183
rl854 n2__i1__net1 n4__i1__net1 56.5719
rl855 i0__net1 n2__i0__net1 56.5719
rl856 n2__i0__net1 n3__i0__net1 48.1183
rl857 n2__i0__net1 n4__i0__net1 56.5719
rl858 n9__i13__net1 n10__i13__net1 87.2876
rl859 n9__i13__net2 n10__i13__net2 87.2876
rl860 i13__i19__i4__net2 n2__i13__i19__i4__net2 82.6365
rl861 i13__i18__i4__net2 n2__i13__i18__i4__net2 82.6365
rl862 n5__i13__net11 n6__i13__net11 56.5719
rl863 n6__i13__net11 n7__i13__net11 48.1183
rl864 n6__i13__net11 n8__i13__net11 56.5719
rl865 n5__i13__net12 n6__i13__net12 56.5719
rl866 n6__i13__net12 n7__i13__net12 48.1183
rl867 n6__i13__net12 n8__i13__net12 56.5719
rl868 n16__ck_buff n17__ck_buff 87.898
rl869 n19__ck_b n20__ck_b 126.36
rl870 n21__ck_b n22__ck_b 126.36
rl871 n18__ck_buff n19__ck_buff 87.898
rl872 n20__ck_buff n21__ck_buff 87.898
rl873 n23__ck_b n24__ck_b 126.36
rl874 i18__net3 n2__i18__net3 26.7741
rl875 n2__i18__net3 n3__i18__net3 29.8991
rl876 n4__i18__net3 n5__i18__net3 26.7741
rl877 n5__i18__net3 n6__i18__net3 29.8991
rl878 n7__i18__net3 n8__i18__net3 26.7741
rl879 n8__i18__net3 n9__i18__net3 29.8991
rl880 i13__net7 n2__i13__net7 137.341
rl881 n2__i13__net7 n3__i13__net7 48.1183
rl882 n2__i13__net7 n4__i13__net7 68.1104
rl883 i13__net17 n2__i13__net17 41.1873
rl884 n2__i13__net17 n3__i13__net17 45
rl885 n2__i13__net17 n4__i13__net17 118.11
rl886 i2__net75 n2__i2__net75 9.7184
rl887 i2__net75 n3__i2__net75 11.2742
rl888 i1__net75 n2__i1__net75 11.2742
rl889 i1__net75 n3__i1__net75 9.7184
rl890 i0__net75 n2__i0__net75 9.7184
rl891 i0__net75 n3__i0__net75 11.2742
rl892 n10__i18__net3 n11__i18__net3 26.7741
rl893 n11__i18__net3 n12__i18__net3 29.8991
rl894 i13__net18 n2__i13__net18 60.4181
rl895 n2__i13__net18 n3__i13__net18 48.1183
rl896 n2__i13__net18 n4__i13__net18 145.033
rl897 i13__net23 n2__i13__net23 98.8796
rl898 n2__i13__net23 n3__i13__net23 45
rl899 n2__i13__net23 n4__i13__net23 60.4181
rl900 n13__i18__net3 n14__i18__net3 26.7741
rl901 n14__i18__net3 n15__i18__net3 29.8991
rl902 n20__reset_buff n21__reset_buff 98.1035
rl903 n22__reset_buff n23__reset_buff 98.1035
rl904 n24__reset_buff n25__reset_buff 98.1035
rl905 i13__i20__net1 n2__i13__i20__net1 56.5719
rl906 n2__i13__i20__net1 n3__i13__i20__net1 48.1183
rl907 n2__i13__i20__net1 n4__i13__i20__net1 56.5719
rl908 i13__net3 n2__i13__net3 49.0903
rl909 n2__i13__net3 n3__i13__net3 49.0903
rl910 n16__i18__net3 n17__i18__net3 26.7741
rl911 n17__i18__net3 n18__i18__net3 29.8991
rl912 i2__net74 n2__i2__net74 56.5719
rl913 n2__i2__net74 n3__i2__net74 23.6889
rl914 n3__i2__net74 n4__i2__net74 50.6296
rl915 n2__i2__net74 n5__i2__net74 56.5719
rl916 n3__i2__net74 n6__i2__net74 55.6157
rl917 n3__i2__net74 n7__i2__net74 55.6157
rl918 i1__net74 n2__i1__net74 56.5719
rl919 n2__i1__net74 n3__i1__net74 23.6889
rl920 n3__i1__net74 n4__i1__net74 50.6296
rl921 n2__i1__net74 n5__i1__net74 56.5719
rl922 n3__i1__net74 n6__i1__net74 55.6157
rl923 n3__i1__net74 n7__i1__net74 55.6157
rl924 i0__net74 n2__i0__net74 56.5719
rl925 n2__i0__net74 n3__i0__net74 23.6889
rl926 n3__i0__net74 n4__i0__net74 50.6296
rl927 n2__i0__net74 n5__i0__net74 56.5719
rl928 n3__i0__net74 n6__i0__net74 55.6157
rl929 n3__i0__net74 n7__i0__net74 55.6157
rl930 n5__i13__net18 n6__i13__net18 56.5719
rl931 n6__i13__net18 n7__i13__net18 48.1183
rl932 n6__i13__net18 n8__i13__net18 56.5719
rl933 n19__i18__net3 n20__i18__net3 26.7741
rl934 n20__i18__net3 n21__i18__net3 29.8991
rl935 n22__i18__net3 n23__i18__net3 26.7741
rl936 n23__i18__net3 n24__i18__net3 29.8991
rl937 n9__i13__net18 n10__i13__net18 87.2876
rl938 n25__ck_b n26__ck_b 87.898
rl939 n28__ck_buff n29__ck_buff 126.36
rl940 n30__ck_buff n31__ck_buff 126.36
rl941 n27__ck_b n28__ck_b 87.898
rl942 n29__ck_b n30__ck_b 87.898
rl943 n32__ck_buff n33__ck_buff 126.36
rl944 i13__i20__i4__net2 n2__i13__i20__i4__net2 82.6365
rl945 n25__i18__net3 n26__i18__net3 26.7741
rl946 n26__i18__net3 n27__i18__net3 29.8991
rl947 n5__i13__net7 n6__i13__net7 56.5719
rl948 n6__i13__net7 n7__i13__net7 48.1183
rl949 n6__i13__net7 n8__i13__net7 56.5719
rl950 n28__i18__net3 n29__i18__net3 26.7741
rl951 n29__i18__net3 n30__i18__net3 29.8991
rl952 n1__serial_out n2__serial_out 59.0671
rl953 i2__net77 n2__i2__net77 9.7184
rl954 i2__net77 n3__i2__net77 11.2742
rl955 i1__net77 n2__i1__net77 11.2742
rl956 i1__net77 n3__i1__net77 9.7184
rl957 i0__net77 n2__i0__net77 9.7184
rl958 i0__net77 n3__i0__net77 11.2742
rl959 n15__reset_b n16__reset_b 74.5009
rl960 n17__reset_b n18__reset_b 74.5009
rl961 n19__reset_b n20__reset_b 74.5009
rl962 n3__serial_out n4__serial_out 59.0671
rl963 n5__serial_out n6__serial_out 59.0671
rl964 i2__net76 n2__i2__net76 56.5719
rl965 n2__i2__net76 n3__i2__net76 23.6889
rl966 n3__i2__net76 n4__i2__net76 50.6296
rl967 n2__i2__net76 n5__i2__net76 56.5719
rl968 n3__i2__net76 n6__i2__net76 55.6157
rl969 n3__i2__net76 n7__i2__net76 55.6157
rl970 i1__net76 n2__i1__net76 56.5719
rl971 n2__i1__net76 n3__i1__net76 23.6889
rl972 n3__i1__net76 n4__i1__net76 50.6296
rl973 n2__i1__net76 n5__i1__net76 56.5719
rl974 n3__i1__net76 n6__i1__net76 55.6157
rl975 n3__i1__net76 n7__i1__net76 55.6157
rl976 i0__net76 n2__i0__net76 56.5719
rl977 n2__i0__net76 n3__i0__net76 23.6889
rl978 n3__i0__net76 n4__i0__net76 50.6296
rl979 n2__i0__net76 n5__i0__net76 56.5719
rl980 n3__i0__net76 n6__i0__net76 55.6157
rl981 n3__i0__net76 n7__i0__net76 55.6157
rl982 i12__bio n2__i12__bio 80.264
rl983 n4__i2__net77 n5__i2__net77 49.0903
rl984 n5__i2__net77 n6__i2__net77 49.0903
rl985 n4__i1__net77 n5__i1__net77 49.0903
rl986 n5__i1__net77 n6__i1__net77 49.0903
rl987 n4__i0__net77 n5__i0__net77 49.0903
rl988 n5__i0__net77 n6__i0__net77 49.0903
rl989 i12__bcore_bar n2__i12__bcore_bar 58.0255
rl990 n7__serial_out n8__serial_out 56.5719
rl991 n8__serial_out n9__serial_out 50.013
rl992 n8__serial_out n10__serial_out 56.5719
rl993 n8__net4 n9__net4 56.5719
rl994 n9__net4 n10__net4 50.013
rl995 n9__net4 n11__net4 56.5719
rl996 n6__net3 n7__net3 56.5719
rl997 n7__net3 n8__net3 50.013
rl998 n7__net3 n9__net3 56.5719
rl999 n3__i12__bcore_bar n4__i12__bcore_bar 58.0255
rl1000 i18__net2 n2__i18__net2 22.3882
rl1001 n2__i18__net2 n3__i18__net2 47.355
rl1002 n3__i18__net2 n4__i18__net2 42.3089
rl1003 n4__i18__net2 n5__i18__net2 36.8896
rl1004 n5__i18__net2 n6__i18__net2 30.5862
rl1005 n2__i18__net2 n7__i18__net2 27.5965
rl1006 n3__i18__net2 n8__i18__net2 30.2243
rl1007 n3__i18__net2 n9__i18__net2 25.0159
rl1008 n4__i18__net2 n10__i18__net2 30.2243
rl1009 n4__i18__net2 n11__i18__net2 25.0159
rl1010 n5__i18__net2 n12__i18__net2 25.3779
rl1011 n5__i12__bcore_bar n6__i12__bcore_bar 58.0255
rl1012 serial_out_b_high n2__serial_out_b_high 59.3399
rl1013 n10__r0 n11__r0 56.5719
rl1014 n11__r0 n12__r0 45
rl1015 n11__r0 n13__r0 56.5719
rl1016 n5__r2 n6__r2 56.5719
rl1017 n6__r2 n7__r2 45
rl1018 n6__r2 n8__r2 56.5719
rl1019 r1 n2__r1 56.5719
rl1020 n2__r1 n3__r1 45
rl1021 n2__r1 n4__r1 56.5719
rl1022 i18__net1 n2__i18__net1 21.3465
rl1023 n2__i18__net1 n3__i18__net1 41.9357
rl1024 n3__i18__net1 n4__i18__net1 30.5862
rl1025 n2__i18__net1 n5__i18__net1 27.5965
rl1026 n3__i18__net1 n6__i18__net1 24.3362
rl1027 n11__serial_out n12__serial_out 58.6166
rl1028 n12__serial_out n13__serial_out 133.617
rl1029 n3__serial_out_b_high n4__serial_out_b_high 17.1921
rl1030 n3__serial_out_b_high n5__serial_out_b_high 16.1505
rl1031 net7 n2__net7 56.5719
rl1032 n2__net7 n3__net7 23.6889
rl1033 n3__net7 n4__net7 26.2002
rl1034 n4__net7 n5__net7 45
rl1035 n2__net7 n6__net7 56.5719
rl1036 n3__net7 n7__net7 55.6157
rl1037 n3__net7 n8__net7 55.6157
rl1038 n4__net7 n9__net7 55.6157
rl1039 n4__net7 n10__net7 55.6157
rl1040 net6 n2__net6 56.5719
rl1041 n2__net6 n3__net6 23.6889
rl1042 n3__net6 n4__net6 26.2002
rl1043 n4__net6 n5__net6 45
rl1044 n2__net6 n6__net6 56.5719
rl1045 n3__net6 n7__net6 55.6157
rl1046 n3__net6 n8__net6 55.6157
rl1047 n4__net6 n9__net6 55.6157
rl1048 n4__net6 n10__net6 55.6157
rl1049 net8 n2__net8 56.5719
rl1050 n2__net8 n3__net8 23.6889
rl1051 n3__net8 n4__net8 26.2002
rl1052 n4__net8 n5__net8 45
rl1053 n2__net8 n6__net8 56.5719
rl1054 n3__net8 n7__net8 55.6157
rl1055 n3__net8 n8__net8 55.6157
rl1056 n4__net8 n9__net8 55.6157
rl1057 n4__net8 n10__net8 55.6157
rl1058 serial_out_b_high_buff n2__serial_out_b_high_buff 21.3465
rl1059 n2__serial_out_b_high_buff n3__serial_out_b_high_buff 27.5965
mi40__m2 n7__serial_out_b_high_buff n5__serial_out_b_high n685__vddio n683__vddio g45p2svt L=150e-9 W=640e-9 AD=96e-15 AS=96e-15 PD=1.58e-6 PS=1.58e-6 NRD=468.75e-3 NRS=468.75e-3 M=1
mi18__m17_99__rcx n35__r_out n18__i18__net5 n952__vddio n686__vddio g45p2svt L=150e-9 W=8.22e-6 AD=1.644e-12 AS=1.644e-12 PD=16.84e-6 PS=16.84e-6 NRD=468.75e-3 NRS=468.75e-3 M=1
mi18__m17_98__rcx n956__vddio n15__i18__net5 n35__r_out n686__vddio g45p2svt L=150e-9 W=8.22e-6 AD=1.644e-12 AS=1.644e-12 PD=16.84e-6 PS=16.84e-6 NRD=468.75e-3 NRS=468.75e-3 M=1
mi18__m17_97__rcx n19__r_out n12__i18__net5 n956__vddio n686__vddio g45p2svt L=150e-9 W=8.22e-6 AD=1.644e-12 AS=1.644e-12 PD=16.84e-6 PS=16.84e-6 NRD=468.75e-3 NRS=468.75e-3 M=1
mi18__m17_96__rcx n960__vddio n9__i18__net5 n19__r_out n686__vddio g45p2svt L=150e-9 W=8.22e-6 AD=1.644e-12 AS=1.644e-12 PD=16.84e-6 PS=16.84e-6 NRD=468.75e-3 NRS=468.75e-3 M=1
mi18__m17_95__rcx n11__r_out n6__i18__net5 n960__vddio n686__vddio g45p2svt L=150e-9 W=8.22e-6 AD=1.644e-12 AS=1.644e-12 PD=16.84e-6 PS=16.84e-6 NRD=468.75e-3 NRS=468.75e-3 M=1
mi18__m17_94__rcx n762__vddio n3__i18__net5 n11__r_out n686__vddio g45p2svt L=150e-9 W=8.22e-6 AD=1.233e-12 AS=1.233e-12 PD=16.79e-6 PS=16.79e-6 NRD=468.75e-3 NRS=468.75e-3 M=1
mi18__m17_93__rcx n76__r_out n36__i18__net5 n940__vddio n686__vddio g45p2svt L=150e-9 W=8.22e-6 AD=1.644e-12 AS=1.644e-12 PD=16.84e-6 PS=16.84e-6 NRD=468.75e-3 NRS=468.75e-3 M=1
mi18__m17_92__rcx n944__vddio n33__i18__net5 n76__r_out n686__vddio g45p2svt L=150e-9 W=8.22e-6 AD=1.644e-12 AS=1.644e-12 PD=16.84e-6 PS=16.84e-6 NRD=468.75e-3 NRS=468.75e-3 M=1
mi18__m17_91__rcx n61__r_out n30__i18__net5 n944__vddio n686__vddio g45p2svt L=150e-9 W=8.22e-6 AD=1.644e-12 AS=1.644e-12 PD=16.84e-6 PS=16.84e-6 NRD=468.75e-3 NRS=468.75e-3 M=1
mi18__m17_90__rcx n948__vddio n27__i18__net5 n61__r_out n686__vddio g45p2svt L=150e-9 W=8.22e-6 AD=1.644e-12 AS=1.644e-12 PD=16.84e-6 PS=16.84e-6 NRD=468.75e-3 NRS=468.75e-3 M=1
mi18__m17_89__rcx n50__r_out n24__i18__net5 n948__vddio n686__vddio g45p2svt L=150e-9 W=8.22e-6 AD=1.644e-12 AS=1.644e-12 PD=16.84e-6 PS=16.84e-6 NRD=468.75e-3 NRS=468.75e-3 M=1
mi18__m17_88__rcx n952__vddio n21__i18__net5 n50__r_out n686__vddio g45p2svt L=150e-9 W=8.22e-6 AD=1.644e-12 AS=1.644e-12 PD=16.84e-6 PS=16.84e-6 NRD=468.75e-3 NRS=468.75e-3 M=1
mi18__m17_87__rcx n940__vddio n39__i18__net5 n84__r_out n686__vddio g45p2svt L=150e-9 W=8.22e-6 AD=1.644e-12 AS=1.644e-12 PD=16.84e-6 PS=16.84e-6 NRD=468.75e-3 NRS=468.75e-3 M=1
mi18__m17_86__rcx n928__vddio n65__i18__net5 n128__r_out n686__vddio g45p2svt L=150e-9 W=8.22e-6 AD=1.644e-12 AS=1.644e-12 PD=16.84e-6 PS=16.84e-6 NRD=468.75e-3 NRS=468.75e-3 M=1
mi18__m17_85__rcx n115__r_out n62__i18__net5 n928__vddio n686__vddio g45p2svt L=150e-9 W=8.22e-6 AD=1.644e-12 AS=1.644e-12 PD=16.84e-6 PS=16.84e-6 NRD=468.75e-3 NRS=468.75e-3 M=1
mi18__m17_84__rcx n932__vddio n55__i18__net5 n115__r_out n686__vddio g45p2svt L=150e-9 W=8.22e-6 AD=1.644e-12 AS=1.644e-12 PD=16.84e-6 PS=16.84e-6 NRD=468.75e-3 NRS=468.75e-3 M=1
mi18__m17_83__rcx n102__r_out n52__i18__net5 n932__vddio n686__vddio g45p2svt L=150e-9 W=8.22e-6 AD=1.644e-12 AS=1.644e-12 PD=16.84e-6 PS=16.84e-6 NRD=468.75e-3 NRS=468.75e-3 M=1
mi18__m17_82__rcx n936__vddio n45__i18__net5 n102__r_out n686__vddio g45p2svt L=150e-9 W=8.22e-6 AD=1.644e-12 AS=1.644e-12 PD=16.84e-6 PS=16.84e-6 NRD=468.75e-3 NRS=468.75e-3 M=1
mi18__m17_81__rcx n84__r_out n42__i18__net5 n936__vddio n686__vddio g45p2svt L=150e-9 W=8.22e-6 AD=1.644e-12 AS=1.644e-12 PD=16.84e-6 PS=16.84e-6 NRD=468.75e-3 NRS=468.75e-3 M=1
mi18__m17_80__rcx n916__vddio n97__i18__net5 n165__r_out n686__vddio g45p2svt L=150e-9 W=8.22e-6 AD=1.644e-12 AS=1.644e-12 PD=16.84e-6 PS=16.84e-6 NRD=468.75e-3 NRS=468.75e-3 M=1
mi18__m17_79__rcx n149__r_out n92__i18__net5 n916__vddio n686__vddio g45p2svt L=150e-9 W=8.22e-6 AD=1.644e-12 AS=1.644e-12 PD=16.84e-6 PS=16.84e-6 NRD=468.75e-3 NRS=468.75e-3 M=1
mi18__m17_78__rcx n920__vddio n87__i18__net5 n149__r_out n686__vddio g45p2svt L=150e-9 W=8.22e-6 AD=1.644e-12 AS=1.644e-12 PD=16.84e-6 PS=16.84e-6 NRD=468.75e-3 NRS=468.75e-3 M=1
mi18__m17_77__rcx n136__r_out n80__i18__net5 n920__vddio n686__vddio g45p2svt L=150e-9 W=8.22e-6 AD=1.644e-12 AS=1.644e-12 PD=16.84e-6 PS=16.84e-6 NRD=468.75e-3 NRS=468.75e-3 M=1
mi18__m17_76__rcx n924__vddio n75__i18__net5 n136__r_out n686__vddio g45p2svt L=150e-9 W=8.22e-6 AD=1.644e-12 AS=1.644e-12 PD=16.84e-6 PS=16.84e-6 NRD=468.75e-3 NRS=468.75e-3 M=1
mi18__m17_75__rcx n128__r_out n70__i18__net5 n924__vddio n686__vddio g45p2svt L=150e-9 W=8.22e-6 AD=1.644e-12 AS=1.644e-12 PD=16.84e-6 PS=16.84e-6 NRD=468.75e-3 NRS=468.75e-3 M=1
mi18__m17_74__rcx n904__vddio n125__i18__net5 n206__r_out n686__vddio g45p2svt L=150e-9 W=8.22e-6 AD=1.644e-12 AS=1.644e-12 PD=16.84e-6 PS=16.84e-6 NRD=468.75e-3 NRS=468.75e-3 M=1
mi18__m17_73__rcx n191__r_out n122__i18__net5 n904__vddio n686__vddio g45p2svt L=150e-9 W=8.22e-6 AD=1.644e-12 AS=1.644e-12 PD=16.84e-6 PS=16.84e-6 NRD=468.75e-3 NRS=468.75e-3 M=1
mi18__m17_72__rcx n908__vddio n117__i18__net5 n191__r_out n686__vddio g45p2svt L=150e-9 W=8.22e-6 AD=1.644e-12 AS=1.644e-12 PD=16.84e-6 PS=16.84e-6 NRD=468.75e-3 NRS=468.75e-3 M=1
mi18__m17_71__rcx n180__r_out n112__i18__net5 n908__vddio n686__vddio g45p2svt L=150e-9 W=8.22e-6 AD=1.644e-12 AS=1.644e-12 PD=16.84e-6 PS=16.84e-6 NRD=468.75e-3 NRS=468.75e-3 M=1
mi18__m17_70__rcx n912__vddio n105__i18__net5 n180__r_out n686__vddio g45p2svt L=150e-9 W=8.22e-6 AD=1.644e-12 AS=1.644e-12 PD=16.84e-6 PS=16.84e-6 NRD=468.75e-3 NRS=468.75e-3 M=1
mi18__m17_69__rcx n165__r_out n102__i18__net5 n912__vddio n686__vddio g45p2svt L=150e-9 W=8.22e-6 AD=1.644e-12 AS=1.644e-12 PD=16.84e-6 PS=16.84e-6 NRD=468.75e-3 NRS=468.75e-3 M=1
mi18__m17_68__rcx n892__vddio n155__i18__net5 n245__r_out n686__vddio g45p2svt L=150e-9 W=8.22e-6 AD=1.644e-12 AS=1.644e-12 PD=16.84e-6 PS=16.84e-6 NRD=468.75e-3 NRS=468.75e-3 M=1
mi18__m17_67__rcx n232__r_out n150__i18__net5 n892__vddio n686__vddio g45p2svt L=150e-9 W=8.22e-6 AD=1.644e-12 AS=1.644e-12 PD=16.84e-6 PS=16.84e-6 NRD=468.75e-3 NRS=468.75e-3 M=1
mi18__m17_66__rcx n896__vddio n145__i18__net5 n232__r_out n686__vddio g45p2svt L=150e-9 W=8.22e-6 AD=1.644e-12 AS=1.644e-12 PD=16.84e-6 PS=16.84e-6 NRD=468.75e-3 NRS=468.75e-3 M=1
mi18__m17_65__rcx n214__r_out n140__i18__net5 n896__vddio n686__vddio g45p2svt L=150e-9 W=8.22e-6 AD=1.644e-12 AS=1.644e-12 PD=16.84e-6 PS=16.84e-6 NRD=468.75e-3 NRS=468.75e-3 M=1
mi18__m17_64__rcx n900__vddio n137__i18__net5 n214__r_out n686__vddio g45p2svt L=150e-9 W=8.22e-6 AD=1.644e-12 AS=1.644e-12 PD=16.84e-6 PS=16.84e-6 NRD=468.75e-3 NRS=468.75e-3 M=1
mi18__m17_63__rcx n206__r_out n131__i18__net5 n900__vddio n686__vddio g45p2svt L=150e-9 W=8.22e-6 AD=1.644e-12 AS=1.644e-12 PD=16.84e-6 PS=16.84e-6 NRD=468.75e-3 NRS=468.75e-3 M=1
mi18__m17_62__rcx n245__r_out n162__i18__net5 n888__vddio n686__vddio g45p2svt L=150e-9 W=8.22e-6 AD=1.644e-12 AS=1.644e-12 PD=16.84e-6 PS=16.84e-6 NRD=468.75e-3 NRS=468.75e-3 M=1
mi18__m17_61__rcx n279__r_out n190__i18__net5 n876__vddio n686__vddio g45p2svt L=150e-9 W=8.22e-6 AD=1.644e-12 AS=1.644e-12 PD=16.84e-6 PS=16.84e-6 NRD=468.75e-3 NRS=468.75e-3 M=1
mi18__m17_60__rcx n880__vddio n187__i18__net5 n279__r_out n686__vddio g45p2svt L=150e-9 W=8.22e-6 AD=1.644e-12 AS=1.644e-12 PD=16.84e-6 PS=16.84e-6 NRD=468.75e-3 NRS=468.75e-3 M=1
mi18__m17_59__rcx n271__r_out n181__i18__net5 n880__vddio n686__vddio g45p2svt L=150e-9 W=8.22e-6 AD=1.644e-12 AS=1.644e-12 PD=16.84e-6 PS=16.84e-6 NRD=468.75e-3 NRS=468.75e-3 M=1
mi18__m17_58__rcx n884__vddio n175__i18__net5 n271__r_out n686__vddio g45p2svt L=150e-9 W=8.22e-6 AD=1.644e-12 AS=1.644e-12 PD=16.84e-6 PS=16.84e-6 NRD=468.75e-3 NRS=468.75e-3 M=1
mi18__m17_57__rcx n258__r_out n172__i18__net5 n884__vddio n686__vddio g45p2svt L=150e-9 W=8.22e-6 AD=1.644e-12 AS=1.644e-12 PD=16.84e-6 PS=16.84e-6 NRD=468.75e-3 NRS=468.75e-3 M=1
mi18__m17_56__rcx n888__vddio n166__i18__net5 n258__r_out n686__vddio g45p2svt L=150e-9 W=8.22e-6 AD=1.644e-12 AS=1.644e-12 PD=16.84e-6 PS=16.84e-6 NRD=468.75e-3 NRS=468.75e-3 M=1
mi18__m17_55__rcx n323__r_out n220__i18__net5 n864__vddio n686__vddio g45p2svt L=150e-9 W=8.22e-6 AD=1.644e-12 AS=1.644e-12 PD=16.84e-6 PS=16.84e-6 NRD=468.75e-3 NRS=468.75e-3 M=1
mi18__m17_54__rcx n868__vddio n216__i18__net5 n323__r_out n686__vddio g45p2svt L=150e-9 W=8.22e-6 AD=1.644e-12 AS=1.644e-12 PD=16.84e-6 PS=16.84e-6 NRD=468.75e-3 NRS=468.75e-3 M=1
mi18__m17_53__rcx n310__r_out n210__i18__net5 n868__vddio n686__vddio g45p2svt L=150e-9 W=8.22e-6 AD=1.644e-12 AS=1.644e-12 PD=16.84e-6 PS=16.84e-6 NRD=468.75e-3 NRS=468.75e-3 M=1
mi18__m17_52__rcx n872__vddio n205__i18__net5 n310__r_out n686__vddio g45p2svt L=150e-9 W=8.22e-6 AD=1.644e-12 AS=1.644e-12 PD=16.84e-6 PS=16.84e-6 NRD=468.75e-3 NRS=468.75e-3 M=1
mi18__m17_51__rcx n297__r_out n201__i18__net5 n872__vddio n686__vddio g45p2svt L=150e-9 W=8.22e-6 AD=1.644e-12 AS=1.644e-12 PD=16.84e-6 PS=16.84e-6 NRD=468.75e-3 NRS=468.75e-3 M=1
mi18__m17_50__rcx n876__vddio n195__i18__net5 n297__r_out n686__vddio g45p2svt L=150e-9 W=8.22e-6 AD=1.644e-12 AS=1.644e-12 PD=16.84e-6 PS=16.84e-6 NRD=468.75e-3 NRS=468.75e-3 M=1
mi18__m17_49__rcx n360__r_out n252__i18__net5 n852__vddio n686__vddio g45p2svt L=150e-9 W=8.22e-6 AD=1.644e-12 AS=1.644e-12 PD=16.84e-6 PS=16.84e-6 NRD=468.75e-3 NRS=468.75e-3 M=1
mi18__m17_48__rcx n856__vddio n247__i18__net5 n360__r_out n686__vddio g45p2svt L=150e-9 W=8.22e-6 AD=1.644e-12 AS=1.644e-12 PD=16.84e-6 PS=16.84e-6 NRD=468.75e-3 NRS=468.75e-3 M=1
mi18__m17_47__rcx n344__r_out n242__i18__net5 n856__vddio n686__vddio g45p2svt L=150e-9 W=8.22e-6 AD=1.644e-12 AS=1.644e-12 PD=16.84e-6 PS=16.84e-6 NRD=468.75e-3 NRS=468.75e-3 M=1
mi18__m17_46__rcx n860__vddio n237__i18__net5 n344__r_out n686__vddio g45p2svt L=150e-9 W=8.22e-6 AD=1.644e-12 AS=1.644e-12 PD=16.84e-6 PS=16.84e-6 NRD=468.75e-3 NRS=468.75e-3 M=1
mi18__m17_45__rcx n336__r_out n230__i18__net5 n860__vddio n686__vddio g45p2svt L=150e-9 W=8.22e-6 AD=1.644e-12 AS=1.644e-12 PD=16.84e-6 PS=16.84e-6 NRD=468.75e-3 NRS=468.75e-3 M=1
mi18__m17_44__rcx n864__vddio n225__i18__net5 n336__r_out n686__vddio g45p2svt L=150e-9 W=8.22e-6 AD=1.644e-12 AS=1.644e-12 PD=16.84e-6 PS=16.84e-6 NRD=468.75e-3 NRS=468.75e-3 M=1
mi18__m17_43__rcx n399__r_out n280__i18__net5 n840__vddio n686__vddio g45p2svt L=150e-9 W=8.22e-6 AD=1.644e-12 AS=1.644e-12 PD=16.84e-6 PS=16.84e-6 NRD=468.75e-3 NRS=468.75e-3 M=1
mi18__m17_42__rcx n844__vddio n277__i18__net5 n399__r_out n686__vddio g45p2svt L=150e-9 W=8.22e-6 AD=1.644e-12 AS=1.644e-12 PD=16.84e-6 PS=16.84e-6 NRD=468.75e-3 NRS=468.75e-3 M=1
mi18__m17_41__rcx n386__r_out n270__i18__net5 n844__vddio n686__vddio g45p2svt L=150e-9 W=8.22e-6 AD=1.644e-12 AS=1.644e-12 PD=16.84e-6 PS=16.84e-6 NRD=468.75e-3 NRS=468.75e-3 M=1
mi18__m17_40__rcx n848__vddio n267__i18__net5 n386__r_out n686__vddio g45p2svt L=150e-9 W=8.22e-6 AD=1.644e-12 AS=1.644e-12 PD=16.84e-6 PS=16.84e-6 NRD=468.75e-3 NRS=468.75e-3 M=1
mi18__m17_39__rcx n375__r_out n260__i18__net5 n848__vddio n686__vddio g45p2svt L=150e-9 W=8.22e-6 AD=1.644e-12 AS=1.644e-12 PD=16.84e-6 PS=16.84e-6 NRD=468.75e-3 NRS=468.75e-3 M=1
mi18__m17_38__rcx n852__vddio n255__i18__net5 n375__r_out n686__vddio g45p2svt L=150e-9 W=8.22e-6 AD=1.644e-12 AS=1.644e-12 PD=16.84e-6 PS=16.84e-6 NRD=468.75e-3 NRS=468.75e-3 M=1
mi18__m17_37__rcx n840__vddio n285__i18__net5 n409__r_out n686__vddio g45p2svt L=150e-9 W=8.22e-6 AD=1.644e-12 AS=1.644e-12 PD=16.84e-6 PS=16.84e-6 NRD=468.75e-3 NRS=468.75e-3 M=1
mi18__m17_36__rcx n828__vddio n315__i18__net5 n450__r_out n686__vddio g45p2svt L=150e-9 W=8.22e-6 AD=1.644e-12 AS=1.644e-12 PD=16.84e-6 PS=16.84e-6 NRD=468.75e-3 NRS=468.75e-3 M=1
mi18__m17_35__rcx n442__r_out n312__i18__net5 n828__vddio n686__vddio g45p2svt L=150e-9 W=8.22e-6 AD=1.644e-12 AS=1.644e-12 PD=16.84e-6 PS=16.84e-6 NRD=468.75e-3 NRS=468.75e-3 M=1
mi18__m17_34__rcx n832__vddio n305__i18__net5 n442__r_out n686__vddio g45p2svt L=150e-9 W=8.22e-6 AD=1.644e-12 AS=1.644e-12 PD=16.84e-6 PS=16.84e-6 NRD=468.75e-3 NRS=468.75e-3 M=1
mi18__m17_33__rcx n422__r_out n300__i18__net5 n832__vddio n686__vddio g45p2svt L=150e-9 W=8.22e-6 AD=1.644e-12 AS=1.644e-12 PD=16.84e-6 PS=16.84e-6 NRD=468.75e-3 NRS=468.75e-3 M=1
mi18__m17_32__rcx n836__vddio n295__i18__net5 n422__r_out n686__vddio g45p2svt L=150e-9 W=8.22e-6 AD=1.644e-12 AS=1.644e-12 PD=16.84e-6 PS=16.84e-6 NRD=468.75e-3 NRS=468.75e-3 M=1
mi18__m17_31__rcx n409__r_out n290__i18__net5 n836__vddio n686__vddio g45p2svt L=150e-9 W=8.22e-6 AD=1.644e-12 AS=1.644e-12 PD=16.84e-6 PS=16.84e-6 NRD=468.75e-3 NRS=468.75e-3 M=1
mi18__m17_30__rcx n816__vddio n347__i18__net5 n497__r_out n686__vddio g45p2svt L=150e-9 W=8.22e-6 AD=1.644e-12 AS=1.644e-12 PD=16.84e-6 PS=16.84e-6 NRD=468.75e-3 NRS=468.75e-3 M=1
mi18__m17_29__rcx n482__r_out n340__i18__net5 n816__vddio n686__vddio g45p2svt L=150e-9 W=8.22e-6 AD=1.644e-12 AS=1.644e-12 PD=16.84e-6 PS=16.84e-6 NRD=468.75e-3 NRS=468.75e-3 M=1
mi18__m17_28__rcx n820__vddio n337__i18__net5 n482__r_out n686__vddio g45p2svt L=150e-9 W=8.22e-6 AD=1.644e-12 AS=1.644e-12 PD=16.84e-6 PS=16.84e-6 NRD=468.75e-3 NRS=468.75e-3 M=1
mi18__m17_27__rcx n466__r_out n330__i18__net5 n820__vddio n686__vddio g45p2svt L=150e-9 W=8.22e-6 AD=1.644e-12 AS=1.644e-12 PD=16.84e-6 PS=16.84e-6 NRD=468.75e-3 NRS=468.75e-3 M=1
mi18__m17_26__rcx n824__vddio n327__i18__net5 n466__r_out n686__vddio g45p2svt L=150e-9 W=8.22e-6 AD=1.644e-12 AS=1.644e-12 PD=16.84e-6 PS=16.84e-6 NRD=468.75e-3 NRS=468.75e-3 M=1
mi18__m17_25__rcx n450__r_out n322__i18__net5 n824__vddio n686__vddio g45p2svt L=150e-9 W=8.22e-6 AD=1.644e-12 AS=1.644e-12 PD=16.84e-6 PS=16.84e-6 NRD=468.75e-3 NRS=468.75e-3 M=1
mi18__m17_24__rcx n804__vddio n377__i18__net5 n531__r_out n686__vddio g45p2svt L=150e-9 W=8.22e-6 AD=1.644e-12 AS=1.644e-12 PD=16.84e-6 PS=16.84e-6 NRD=468.75e-3 NRS=468.75e-3 M=1
mi18__m17_23__rcx n521__r_out n370__i18__net5 n804__vddio n686__vddio g45p2svt L=150e-9 W=8.22e-6 AD=1.644e-12 AS=1.644e-12 PD=16.84e-6 PS=16.84e-6 NRD=468.75e-3 NRS=468.75e-3 M=1
mi18__m17_22__rcx n808__vddio n367__i18__net5 n521__r_out n686__vddio g45p2svt L=150e-9 W=8.22e-6 AD=1.644e-12 AS=1.644e-12 PD=16.84e-6 PS=16.84e-6 NRD=468.75e-3 NRS=468.75e-3 M=1
mi18__m17_21__rcx n510__r_out n362__i18__net5 n808__vddio n686__vddio g45p2svt L=150e-9 W=8.22e-6 AD=1.644e-12 AS=1.644e-12 PD=16.84e-6 PS=16.84e-6 NRD=468.75e-3 NRS=468.75e-3 M=1
mi18__m17_20__rcx n812__vddio n357__i18__net5 n510__r_out n686__vddio g45p2svt L=150e-9 W=8.22e-6 AD=1.644e-12 AS=1.644e-12 PD=16.84e-6 PS=16.84e-6 NRD=468.75e-3 NRS=468.75e-3 M=1
mi18__m17_19__rcx n497__r_out n350__i18__net5 n812__vddio n686__vddio g45p2svt L=150e-9 W=8.22e-6 AD=1.644e-12 AS=1.644e-12 PD=16.84e-6 PS=16.84e-6 NRD=468.75e-3 NRS=468.75e-3 M=1
mi18__m17_18__rcx n792__vddio n407__i18__net5 n570__r_out n686__vddio g45p2svt L=150e-9 W=8.22e-6 AD=1.644e-12 AS=1.644e-12 PD=16.84e-6 PS=16.84e-6 NRD=468.75e-3 NRS=468.75e-3 M=1
mi18__m17_17__rcx n557__r_out n400__i18__net5 n792__vddio n686__vddio g45p2svt L=150e-9 W=8.22e-6 AD=1.644e-12 AS=1.644e-12 PD=16.84e-6 PS=16.84e-6 NRD=468.75e-3 NRS=468.75e-3 M=1
mi18__m17_16__rcx n796__vddio n397__i18__net5 n557__r_out n686__vddio g45p2svt L=150e-9 W=8.22e-6 AD=1.644e-12 AS=1.644e-12 PD=16.84e-6 PS=16.84e-6 NRD=468.75e-3 NRS=468.75e-3 M=1
mi18__m17_15__rcx n544__r_out n392__i18__net5 n796__vddio n686__vddio g45p2svt L=150e-9 W=8.22e-6 AD=1.644e-12 AS=1.644e-12 PD=16.84e-6 PS=16.84e-6 NRD=468.75e-3 NRS=468.75e-3 M=1
mi18__m17_14__rcx n800__vddio n387__i18__net5 n544__r_out n686__vddio g45p2svt L=150e-9 W=8.22e-6 AD=1.644e-12 AS=1.644e-12 PD=16.84e-6 PS=16.84e-6 NRD=468.75e-3 NRS=468.75e-3 M=1
mi18__m17_13__rcx n531__r_out n380__i18__net5 n800__vddio n686__vddio g45p2svt L=150e-9 W=8.22e-6 AD=1.644e-12 AS=1.644e-12 PD=16.84e-6 PS=16.84e-6 NRD=468.75e-3 NRS=468.75e-3 M=1
mi18__m17_12__rcx n570__r_out n410__i18__net5 n788__vddio n686__vddio g45p2svt L=150e-9 W=8.22e-6 AD=1.644e-12 AS=1.644e-12 PD=16.84e-6 PS=16.84e-6 NRD=468.75e-3 NRS=468.75e-3 M=1
mi18__m17_11__rcx n609__r_out n442__i18__net5 n776__vddio n686__vddio g45p2svt L=150e-9 W=8.22e-6 AD=1.644e-12 AS=1.644e-12 PD=16.84e-6 PS=16.84e-6 NRD=468.75e-3 NRS=468.75e-3 M=1
mi18__m17_10__rcx n780__vddio n437__i18__net5 n609__r_out n686__vddio g45p2svt L=150e-9 W=8.22e-6 AD=1.644e-12 AS=1.644e-12 PD=16.84e-6 PS=16.84e-6 NRD=468.75e-3 NRS=468.75e-3 M=1
mi18__m17_9__rcx n596__r_out n430__i18__net5 n780__vddio n686__vddio g45p2svt L=150e-9 W=8.22e-6 AD=1.644e-12 AS=1.644e-12 PD=16.84e-6 PS=16.84e-6 NRD=468.75e-3 NRS=468.75e-3 M=1
mi18__m17_8__rcx n784__vddio n425__i18__net5 n596__r_out n686__vddio g45p2svt L=150e-9 W=8.22e-6 AD=1.644e-12 AS=1.644e-12 PD=16.84e-6 PS=16.84e-6 NRD=468.75e-3 NRS=468.75e-3 M=1
mi18__m17_7__rcx n583__r_out n421__i18__net5 n784__vddio n686__vddio g45p2svt L=150e-9 W=8.22e-6 AD=1.644e-12 AS=1.644e-12 PD=16.84e-6 PS=16.84e-6 NRD=468.75e-3 NRS=468.75e-3 M=1
mi18__m17_6__rcx n788__vddio n415__i18__net5 n583__r_out n686__vddio g45p2svt L=150e-9 W=8.22e-6 AD=1.644e-12 AS=1.644e-12 PD=16.84e-6 PS=16.84e-6 NRD=468.75e-3 NRS=468.75e-3 M=1
mi18__m17_5__rcx n768__vddio n465__i18__net5 n648__r_out n686__vddio g45p2svt L=150e-9 W=8.22e-6 AD=1.644e-12 AS=1.644e-12 PD=16.84e-6 PS=16.84e-6 NRD=468.75e-3 NRS=468.75e-3 M=1
mi18__m17_4__rcx n635__r_out n460__i18__net5 n768__vddio n686__vddio g45p2svt L=150e-9 W=8.22e-6 AD=1.644e-12 AS=1.644e-12 PD=16.84e-6 PS=16.84e-6 NRD=468.75e-3 NRS=468.75e-3 M=1
mi18__m17_3__rcx n772__vddio n455__i18__net5 n635__r_out n686__vddio g45p2svt L=150e-9 W=8.22e-6 AD=1.644e-12 AS=1.644e-12 PD=16.84e-6 PS=16.84e-6 NRD=468.75e-3 NRS=468.75e-3 M=1
mi18__m17_2__rcx n622__r_out n452__i18__net5 n772__vddio n686__vddio g45p2svt L=150e-9 W=8.22e-6 AD=1.644e-12 AS=1.644e-12 PD=16.84e-6 PS=16.84e-6 NRD=468.75e-3 NRS=468.75e-3 M=1
mi18__m17_1__rcx n776__vddio n445__i18__net5 n622__r_out n686__vddio g45p2svt L=150e-9 W=8.22e-6 AD=1.644e-12 AS=1.644e-12 PD=16.84e-6 PS=16.84e-6 NRD=468.75e-3 NRS=468.75e-3 M=1
mi18__m17 n648__r_out n472__i18__net5 n699__vddio n686__vddio g45p2svt L=150e-9 W=8.22e-6 AD=1.644e-12 AS=1.644e-12 PD=16.79e-6 PS=16.79e-6 NRD=468.75e-3 NRS=468.75e-3 M=1
mi18__m16_29__rcx n598__vddio n21__i18__net4 n546__i18__net5 n686__vddio g45p2svt L=150e-9 W=7.65e-6 AD=1.53e-12 AS=1.53e-12 PD=15.7e-6 PS=15.7e-6 NRD=468.75e-3 NRS=468.75e-3 M=1
mi18__m16_28__rcx n533__i18__net5 n18__i18__net4 n598__vddio n686__vddio g45p2svt L=150e-9 W=7.65e-6 AD=1.53e-12 AS=1.53e-12 PD=15.7e-6 PS=15.7e-6 NRD=468.75e-3 NRS=468.75e-3 M=1
mi18__m16_27__rcx n602__vddio n15__i18__net4 n533__i18__net5 n686__vddio g45p2svt L=150e-9 W=7.65e-6 AD=1.53e-12 AS=1.53e-12 PD=15.7e-6 PS=15.7e-6 NRD=468.75e-3 NRS=468.75e-3 M=1
mi18__m16_26__rcx n520__i18__net5 n12__i18__net4 n602__vddio n686__vddio g45p2svt L=150e-9 W=7.65e-6 AD=1.53e-12 AS=1.53e-12 PD=15.7e-6 PS=15.7e-6 NRD=468.75e-3 NRS=468.75e-3 M=1
mi18__m16_25__rcx n606__vddio n9__i18__net4 n520__i18__net5 n686__vddio g45p2svt L=150e-9 W=7.65e-6 AD=1.53e-12 AS=1.53e-12 PD=15.7e-6 PS=15.7e-6 NRD=468.75e-3 NRS=468.75e-3 M=1
mi18__m16_24__rcx n510__i18__net5 n6__i18__net4 n606__vddio n686__vddio g45p2svt L=150e-9 W=7.65e-6 AD=1.53e-12 AS=1.53e-12 PD=15.7e-6 PS=15.7e-6 NRD=468.75e-3 NRS=468.75e-3 M=1
mi18__m16_23__rcx n610__vddio n3__i18__net4 n510__i18__net5 n686__vddio g45p2svt L=150e-9 W=7.65e-6 AD=1.1475e-12 AS=1.1475e-12 PD=15.65e-6 PS=15.65e-6 NRD=468.75e-3 NRS=468.75e-3 M=1
mi18__m16_22__rcx n585__i18__net5 n42__i18__net4 n614__vddio n686__vddio g45p2svt L=150e-9 W=7.65e-6 AD=1.53e-12 AS=1.53e-12 PD=15.7e-6 PS=15.7e-6 NRD=468.75e-3 NRS=468.75e-3 M=1
mi18__m16_21__rcx n617__vddio n39__i18__net4 n585__i18__net5 n686__vddio g45p2svt L=150e-9 W=7.65e-6 AD=1.53e-12 AS=1.53e-12 PD=15.7e-6 PS=15.7e-6 NRD=468.75e-3 NRS=468.75e-3 M=1
mi18__m16_20__rcx n572__i18__net5 n36__i18__net4 n617__vddio n686__vddio g45p2svt L=150e-9 W=7.65e-6 AD=1.53e-12 AS=1.53e-12 PD=15.7e-6 PS=15.7e-6 NRD=468.75e-3 NRS=468.75e-3 M=1
mi18__m16_19__rcx n590__vddio n33__i18__net4 n572__i18__net5 n686__vddio g45p2svt L=150e-9 W=7.65e-6 AD=1.53e-12 AS=1.53e-12 PD=15.7e-6 PS=15.7e-6 NRD=468.75e-3 NRS=468.75e-3 M=1
mi18__m16_18__rcx n564__i18__net5 n30__i18__net4 n590__vddio n686__vddio g45p2svt L=150e-9 W=7.65e-6 AD=1.53e-12 AS=1.53e-12 PD=15.7e-6 PS=15.7e-6 NRD=468.75e-3 NRS=468.75e-3 M=1
mi18__m16_17__rcx n594__vddio n27__i18__net4 n564__i18__net5 n686__vddio g45p2svt L=150e-9 W=7.65e-6 AD=1.53e-12 AS=1.53e-12 PD=15.7e-6 PS=15.7e-6 NRD=468.75e-3 NRS=468.75e-3 M=1
mi18__m16_16__rcx n546__i18__net5 n24__i18__net4 n594__vddio n686__vddio g45p2svt L=150e-9 W=7.65e-6 AD=1.53e-12 AS=1.53e-12 PD=15.7e-6 PS=15.7e-6 NRD=468.75e-3 NRS=468.75e-3 M=1
mi18__m16_15__rcx n614__vddio n47__i18__net4 n603__i18__net5 n686__vddio g45p2svt L=150e-9 W=7.65e-6 AD=1.53e-12 AS=1.53e-12 PD=15.7e-6 PS=15.7e-6 NRD=468.75e-3 NRS=468.75e-3 M=1
mi18__m16_14__rcx n642__i18__net5 n82__i18__net4 n572__vddio n686__vddio g45p2svt L=150e-9 W=7.65e-6 AD=1.53e-12 AS=1.53e-12 PD=15.7e-6 PS=15.7e-6 NRD=468.75e-3 NRS=468.75e-3 M=1
mi18__m16_13__rcx n576__vddio n75__i18__net4 n642__i18__net5 n686__vddio g45p2svt L=150e-9 W=7.65e-6 AD=1.53e-12 AS=1.53e-12 PD=15.7e-6 PS=15.7e-6 NRD=468.75e-3 NRS=468.75e-3 M=1
mi18__m16_12__rcx n624__i18__net5 n70__i18__net4 n576__vddio n686__vddio g45p2svt L=150e-9 W=7.65e-6 AD=1.53e-12 AS=1.53e-12 PD=15.7e-6 PS=15.7e-6 NRD=468.75e-3 NRS=468.75e-3 M=1
mi18__m16_11__rcx n580__vddio n65__i18__net4 n624__i18__net5 n686__vddio g45p2svt L=150e-9 W=7.65e-6 AD=1.53e-12 AS=1.53e-12 PD=15.7e-6 PS=15.7e-6 NRD=468.75e-3 NRS=468.75e-3 M=1
mi18__m16_10__rcx n611__i18__net5 n61__i18__net4 n580__vddio n686__vddio g45p2svt L=150e-9 W=7.65e-6 AD=1.53e-12 AS=1.53e-12 PD=15.7e-6 PS=15.7e-6 NRD=468.75e-3 NRS=468.75e-3 M=1
mi18__m16_9__rcx n584__vddio n55__i18__net4 n611__i18__net5 n686__vddio g45p2svt L=150e-9 W=7.65e-6 AD=1.53e-12 AS=1.53e-12 PD=15.7e-6 PS=15.7e-6 NRD=468.75e-3 NRS=468.75e-3 M=1
mi18__m16_8__rcx n603__i18__net5 n50__i18__net4 n584__vddio n686__vddio g45p2svt L=150e-9 W=7.65e-6 AD=1.53e-12 AS=1.53e-12 PD=15.7e-6 PS=15.7e-6 NRD=468.75e-3 NRS=468.75e-3 M=1
mi18__m16_7__rcx n560__vddio n115__i18__net4 n689__i18__net5 n686__vddio g45p2svt L=150e-9 W=7.65e-6 AD=1.53e-12 AS=1.53e-12 PD=15.7e-6 PS=15.7e-6 NRD=468.75e-3 NRS=468.75e-3 M=1
mi18__m16_6__rcx n681__i18__net5 n112__i18__net4 n560__vddio n686__vddio g45p2svt L=150e-9 W=7.65e-6 AD=1.53e-12 AS=1.53e-12 PD=15.7e-6 PS=15.7e-6 NRD=468.75e-3 NRS=468.75e-3 M=1
mi18__m16_5__rcx n564__vddio n105__i18__net4 n681__i18__net5 n686__vddio g45p2svt L=150e-9 W=7.65e-6 AD=1.53e-12 AS=1.53e-12 PD=15.7e-6 PS=15.7e-6 NRD=468.75e-3 NRS=468.75e-3 M=1
mi18__m16_4__rcx n663__i18__net5 n102__i18__net4 n564__vddio n686__vddio g45p2svt L=150e-9 W=7.65e-6 AD=1.53e-12 AS=1.53e-12 PD=15.7e-6 PS=15.7e-6 NRD=468.75e-3 NRS=468.75e-3 M=1
mi18__m16_3__rcx n568__vddio n97__i18__net4 n663__i18__net5 n686__vddio g45p2svt L=150e-9 W=7.65e-6 AD=1.53e-12 AS=1.53e-12 PD=15.7e-6 PS=15.7e-6 NRD=468.75e-3 NRS=468.75e-3 M=1
mi18__m16_2__rcx n650__i18__net5 n90__i18__net4 n568__vddio n686__vddio g45p2svt L=150e-9 W=7.65e-6 AD=1.53e-12 AS=1.53e-12 PD=15.7e-6 PS=15.7e-6 NRD=468.75e-3 NRS=468.75e-3 M=1
mi18__m16_1__rcx n572__vddio n85__i18__net4 n650__i18__net5 n686__vddio g45p2svt L=150e-9 W=7.65e-6 AD=1.53e-12 AS=1.53e-12 PD=15.7e-6 PS=15.7e-6 NRD=468.75e-3 NRS=468.75e-3 M=1
mi18__m9_9__rcx n200__i18__net4 n30__i18__net3 n636__vddio n686__vddio g45p2svt L=150e-9 W=6.28e-6 AD=1.256e-12 AS=1.256e-12 PD=12.91e-6 PS=12.91e-6 NRD=468.75e-3 NRS=468.75e-3 M=1
mi18__m9_8__rcx n643__vddio n27__i18__net3 n200__i18__net4 n686__vddio g45p2svt L=150e-9 W=6.28e-6 AD=1.256e-12 AS=1.256e-12 PD=12.96e-6 PS=12.96e-6 NRD=468.75e-3 NRS=468.75e-3 M=1
mi18__m9_7__rcx n189__i18__net4 n24__i18__net3 n643__vddio n686__vddio g45p2svt L=150e-9 W=6.28e-6 AD=1.256e-12 AS=1.256e-12 PD=12.96e-6 PS=12.96e-6 NRD=468.75e-3 NRS=468.75e-3 M=1
mi18__m9_6__rcx n646__vddio n21__i18__net3 n189__i18__net4 n686__vddio g45p2svt L=150e-9 W=6.28e-6 AD=1.256e-12 AS=1.256e-12 PD=12.96e-6 PS=12.96e-6 NRD=468.75e-3 NRS=468.75e-3 M=1
mi18__m9_5__rcx n183__i18__net4 n18__i18__net3 n646__vddio n686__vddio g45p2svt L=150e-9 W=6.28e-6 AD=1.256e-12 AS=1.256e-12 PD=12.96e-6 PS=12.96e-6 NRD=468.75e-3 NRS=468.75e-3 M=1
mi18__m9_4__rcx n653__vddio n15__i18__net3 n183__i18__net4 n686__vddio g45p2svt L=150e-9 W=6.28e-6 AD=1.256e-12 AS=1.256e-12 PD=12.96e-6 PS=12.96e-6 NRD=468.75e-3 NRS=468.75e-3 M=1
mi18__m9_3__rcx n167__i18__net4 n12__i18__net3 n653__vddio n686__vddio g45p2svt L=150e-9 W=6.28e-6 AD=1.256e-12 AS=1.256e-12 PD=12.96e-6 PS=12.96e-6 NRD=468.75e-3 NRS=468.75e-3 M=1
mi18__m9_2__rcx n656__vddio n9__i18__net3 n167__i18__net4 n686__vddio g45p2svt L=150e-9 W=6.28e-6 AD=1.256e-12 AS=1.256e-12 PD=12.96e-6 PS=12.96e-6 NRD=468.75e-3 NRS=468.75e-3 M=1
mi18__m9_1__rcx n156__i18__net4 n6__i18__net3 n656__vddio n686__vddio g45p2svt L=150e-9 W=6.28e-6 AD=1.256e-12 AS=1.256e-12 PD=12.96e-6 PS=12.96e-6 NRD=468.75e-3 NRS=468.75e-3 M=1
mi18__m9 n650__vddio n3__i18__net3 n156__i18__net4 n686__vddio g45p2svt L=150e-9 W=6.28e-6 AD=942e-15 AS=942e-15 PD=12.91e-6 PS=12.91e-6 NRD=468.75e-3 NRS=468.75e-3 M=1
mi18__m16 n689__i18__net5 n122__i18__net4 n535__vddio n686__vddio g45p2svt L=150e-9 W=7.65e-6 AD=1.53e-12 AS=1.53e-12 PD=15.65e-6 PS=15.65e-6 NRD=468.75e-3 NRS=468.75e-3 M=1
mi18__m6 n9__i18__net1 n3__serial_out_b_high_buff n678__vddio n686__vddio g45p2svt L=150e-9 W=1.32e-6 AD=198e-15 AS=198e-15 PD=2.94e-6 PS=2.94e-6 NRD=468.75e-3 NRS=468.75e-3 M=1
mi18__m7_1__rcx n15__i18__net2 n5__i18__net1 n682__vddio n686__vddio g45p2svt L=150e-9 W=2.38e-6 AD=476e-15 AS=476e-15 PD=5.11e-6 PS=5.11e-6 NRD=468.75e-3 NRS=468.75e-3 M=1
mi18__m7 n681__vddio n4__i18__net1 n15__i18__net2 n686__vddio g45p2svt L=150e-9 W=2.38e-6 AD=357e-15 AS=357e-15 PD=5.11e-6 PS=5.11e-6 NRD=468.75e-3 NRS=468.75e-3 M=1
mi18__m8_3__rcx n56__i18__net3 n7__i18__net2 n659__vddio n686__vddio g45p2svt L=150e-9 W=4.33e-6 AD=866e-15 AS=866e-15 PD=9.01e-6 PS=9.01e-6 NRD=468.75e-3 NRS=468.75e-3 M=1
mi18__m8_2__rcx n664__vddio n8__i18__net2 n56__i18__net3 n686__vddio g45p2svt L=150e-9 W=4.33e-6 AD=866e-15 AS=866e-15 PD=9.06e-6 PS=9.06e-6 NRD=468.75e-3 NRS=468.75e-3 M=1
mi18__m8_1__rcx n58__i18__net3 n10__i18__net2 n664__vddio n686__vddio g45p2svt L=150e-9 W=4.33e-6 AD=866e-15 AS=866e-15 PD=9.06e-6 PS=9.06e-6 NRD=468.75e-3 NRS=468.75e-3 M=1
mi18__m8 n662__vddio n6__i18__net2 n58__i18__net3 n686__vddio g45p2svt L=150e-9 W=4.33e-6 AD=649.5e-15 AS=649.5e-15 PD=9.01e-6 PS=9.01e-6 NRD=468.75e-3 NRS=468.75e-3 M=1
mi12__m0 n5__i12__bio n2__serial_out_b_high n676__vddio n672__vddio g45p2svt L=150e-9 W=320e-9 AD=48e-15 AS=48e-15 PD=939.999e-9 PS=939.999e-9 NRD=468.75e-3 NRS=468.75e-3 M=1
mi12__m1 n6__serial_out_b_high n2__i12__bio n677__vddio n672__vddio g45p2svt L=150e-9 W=320e-9 AD=48e-15 AS=48e-15 PD=939.999e-9 PS=939.999e-9 NRD=468.75e-3 NRS=468.75e-3 M=1
mi36__m2_2__rcx n15__ck_buff n7__net13 n230__vdd n134__vdd g45p1svt L=45e-9 W=480e-9 AD=76.8e-15 AS=76.8e-15 PD=1.26e-6 PS=1.26e-6 NRD=1.16667 NRS=1.16667 M=1
mi36__m2_1__rcx n228__vdd n5__net13 n15__ck_buff n134__vdd g45p1svt L=45e-9 W=480e-9 AD=76.8e-15 AS=76.8e-15 PD=1.28e-6 PS=1.28e-6 NRD=1.16667 NRS=1.16667 M=1
mi36__m2 n26__ck_buff n3__net13 n228__vdd n134__vdd g45p1svt L=45e-9 W=480e-9 AD=67.2e-15 AS=67.2e-15 PD=1.26e-6 PS=1.26e-6 NRD=1.16667 NRS=1.16667 M=1
mi32__m2_2__rcx n11__ck_b n5__net11 n242__vdd n134__vdd g45p1svt L=45e-9 W=480e-9 AD=76.8e-15 AS=76.8e-15 PD=1.26e-6 PS=1.26e-6 NRD=1.16667 NRS=1.16667 M=1
mi32__m2_1__rcx n243__vdd n7__net11 n11__ck_b n134__vdd g45p1svt L=45e-9 W=480e-9 AD=76.8e-15 AS=76.8e-15 PD=1.28e-6 PS=1.28e-6 NRD=1.16667 NRS=1.16667 M=1
mi32__m2 n7__ck_b n9__net11 n243__vdd n134__vdd g45p1svt L=45e-9 W=480e-9 AD=67.2e-15 AS=67.2e-15 PD=1.26e-6 PS=1.26e-6 NRD=1.16667 NRS=1.16667 M=1
mi37__m2_2__rcx n12__reset_buff n7__net14 n377__vdd n293__vdd g45p1svt L=45e-9 W=480e-9 AD=76.8e-15 AS=76.8e-15 PD=1.26e-6 PS=1.26e-6 NRD=1.16667 NRS=1.16667 M=1
mi37__m2_1__rcx n376__vdd n5__net14 n12__reset_buff n293__vdd g45p1svt L=45e-9 W=480e-9 AD=76.8e-15 AS=76.8e-15 PD=1.28e-6 PS=1.28e-6 NRD=1.16667 NRS=1.16667 M=1
mi37__m2 n15__reset_buff n3__net14 n376__vdd n293__vdd g45p1svt L=45e-9 W=480e-9 AD=67.2e-15 AS=67.2e-15 PD=1.26e-6 PS=1.26e-6 NRD=1.16667 NRS=1.16667 M=1
mi33__m2_2__rcx n12__reset_b n5__net12 n382__vdd n293__vdd g45p1svt L=45e-9 W=480e-9 AD=76.8e-15 AS=76.8e-15 PD=1.26e-6 PS=1.26e-6 NRD=1.16667 NRS=1.16667 M=1
mi33__m2_1__rcx n383__vdd n7__net12 n12__reset_b n293__vdd g45p1svt L=45e-9 W=480e-9 AD=76.8e-15 AS=76.8e-15 PD=1.28e-6 PS=1.28e-6 NRD=1.16667 NRS=1.16667 M=1
mi33__m2 n9__reset_b n9__net12 n383__vdd n293__vdd g45p1svt L=45e-9 W=480e-9 AD=67.2e-15 AS=67.2e-15 PD=1.26e-6 PS=1.26e-6 NRD=1.16667 NRS=1.16667 M=1
mi30__m2_2__rcx n16__net11 n6__net9 n239__vdd n134__vdd g45p1svt L=45e-9 W=240e-9 AD=38.4e-15 AS=38.4e-15 PD=780e-9 PS=780e-9 NRD=1.16667 NRS=1.16667 M=1
mi30__m2_1__rcx n240__vdd n8__net9 n16__net11 n134__vdd g45p1svt L=45e-9 W=240e-9 AD=38.4e-15 AS=38.4e-15 PD=800e-9 PS=800e-9 NRD=1.16667 NRS=1.16667 M=1
mi30__m2 n17__net11 n5__net9 n240__vdd n134__vdd g45p1svt L=45e-9 W=240e-9 AD=33.6e-15 AS=33.6e-15 PD=780e-9 PS=780e-9 NRD=1.16667 NRS=1.16667 M=1
mi29__m2_2__rcx n14__r2_buff n9__net6 n351__vdd n293__vdd g45p1svt L=45e-9 W=240e-9 AD=38.4e-15 AS=38.4e-15 PD=780e-9 PS=780e-9 NRD=1.16667 NRS=1.16667 M=1
mi29__m2_1__rcx n291__vdd n7__net6 n14__r2_buff n293__vdd g45p1svt L=45e-9 W=240e-9 AD=38.4e-15 AS=38.4e-15 PD=800e-9 PS=800e-9 NRD=1.16667 NRS=1.16667 M=1
mi29__m2 n8__r2_buff n6__net6 n291__vdd n293__vdd g45p1svt L=45e-9 W=240e-9 AD=33.6e-15 AS=33.6e-15 PD=780e-9 PS=780e-9 NRD=1.16667 NRS=1.16667 M=1
mi31__m2_2__rcx n16__net12 n6__net10 n380__vdd n293__vdd g45p1svt L=45e-9 W=240e-9 AD=38.4e-15 AS=38.4e-15 PD=780e-9 PS=780e-9 NRD=1.16667 NRS=1.16667 M=1
mi31__m2_1__rcx n381__vdd n8__net10 n16__net12 n293__vdd g45p1svt L=45e-9 W=240e-9 AD=38.4e-15 AS=38.4e-15 PD=800e-9 PS=800e-9 NRD=1.16667 NRS=1.16667 M=1
mi31__m2 n17__net12 n5__net10 n381__vdd n293__vdd g45p1svt L=45e-9 W=240e-9 AD=33.6e-15 AS=33.6e-15 PD=780e-9 PS=780e-9 NRD=1.16667 NRS=1.16667 M=1
mi27__m2_2__rcx n14__r0_buff n10__net7 n211__vdd n134__vdd g45p1svt L=45e-9 W=240e-9 AD=38.4e-15 AS=38.4e-15 PD=780e-9 PS=780e-9 NRD=1.16667 NRS=1.16667 M=1
mi27__m2_1__rcx n133__vdd n8__net7 n14__r0_buff n134__vdd g45p1svt L=45e-9 W=240e-9 AD=38.4e-15 AS=38.4e-15 PD=800e-9 PS=800e-9 NRD=1.16667 NRS=1.16667 M=1
mi27__m2 n8__r0_buff net7 n133__vdd n134__vdd g45p1svt L=45e-9 W=240e-9 AD=33.6e-15 AS=33.6e-15 PD=780e-9 PS=780e-9 NRD=1.16667 NRS=1.16667 M=1
mi28__m2_2__rcx n14__r1_buff n10__net8 n350__vdd n293__vdd g45p1svt L=45e-9 W=240e-9 AD=38.4e-15 AS=38.4e-15 PD=780e-9 PS=780e-9 NRD=1.16667 NRS=1.16667 M=1
mi28__m2_1__rcx n349__vdd n8__net8 n14__r1_buff n293__vdd g45p1svt L=45e-9 W=240e-9 AD=38.4e-15 AS=38.4e-15 PD=800e-9 PS=800e-9 NRD=1.16667 NRS=1.16667 M=1
mi28__m2 n8__r1_buff net8 n349__vdd n293__vdd g45p1svt L=45e-9 W=240e-9 AD=33.6e-15 AS=33.6e-15 PD=780e-9 PS=780e-9 NRD=1.16667 NRS=1.16667 M=1
mi34__m2 n13__net13 n29__ck n232__vdd n134__vdd g45p1svt L=45e-9 W=240e-9 AD=33.6e-15 AS=33.6e-15 PD=760e-9 PS=760e-9 NRD=1.16667 NRS=1.16667 M=1
mi16__m2 n13__net9 n24__ck n237__vdd n134__vdd g45p1svt L=45e-9 W=240e-9 AD=33.6e-15 AS=33.6e-15 PD=760e-9 PS=760e-9 NRD=1.16667 NRS=1.16667 M=1
mi23__m2 n12__net6 n8__r2 n353__vdd n293__vdd g45p1svt L=45e-9 W=240e-9 AD=33.6e-15 AS=33.6e-15 PD=760e-9 PS=760e-9 NRD=1.16667 NRS=1.16667 M=1
mi17__m2 n13__net10 n53__reset n379__vdd n293__vdd g45p1svt L=45e-9 W=240e-9 AD=33.6e-15 AS=33.6e-15 PD=760e-9 PS=760e-9 NRD=1.16667 NRS=1.16667 M=1
mi35__m2 n13__net14 n58__reset n378__vdd n293__vdd g45p1svt L=45e-9 W=240e-9 AD=33.6e-15 AS=33.6e-15 PD=760e-9 PS=760e-9 NRD=1.16667 NRS=1.16667 M=1
mi19__m2 n13__net7 n10__r0 n212__vdd n134__vdd g45p1svt L=45e-9 W=240e-9 AD=33.6e-15 AS=33.6e-15 PD=760e-9 PS=760e-9 NRD=1.16667 NRS=1.16667 M=1
mi22__m2 n13__net8 r1 n352__vdd n293__vdd g45p1svt L=45e-9 W=240e-9 AD=33.6e-15 AS=33.6e-15 PD=760e-9 PS=760e-9 NRD=1.16667 NRS=1.16667 M=1
mi2__pm1_1__rcx n11__i2__net75 n7__i2__net74 n220__vdd n134__vdd g45p1svt L=45e-9 W=480e-9 AD=76.8e-15 AS=76.8e-15 PD=1.26e-6 PS=1.26e-6 NRD=1.16667 NRS=1.16667 M=1
mi2__pm1 n219__vdd i2__net74 n11__i2__net75 n134__vdd g45p1svt L=45e-9 W=480e-9 AD=67.2e-15 AS=67.2e-15 PD=1.26e-6 PS=1.26e-6 NRD=1.16667 NRS=1.16667 M=1
mi2__pm8 n13__i2__net76 n26__ck_b n6__i2__net75 n134__vdd g45p1svt L=45e-9 W=120e-9 AD=16.8e-15 AS=16.8e-15 PD=520e-9 PS=520e-9 NRD=1.16667 NRS=1.16667 M=1
mi2__pm10 n218__vdd n3__i2__net77 n9__i2__net76 n134__vdd g45p1svt L=180e-9 W=120e-9 AD=16.8e-15 AS=16.8e-15 PD=520e-9 PS=520e-9 NRD=1.16667 NRS=1.16667 M=1
mi2__pm15 n15__i2__net76 n15__reset_b n217__vdd n134__vdd g45p1svt L=45e-9 W=120e-9 AD=16.8e-15 AS=16.8e-15 PD=520e-9 PS=520e-9 NRD=1.16667 NRS=1.16667 M=1
mi2__pm9_1__rcx n10__i2__net77 n7__i2__net76 n216__vdd n134__vdd g45p1svt L=45e-9 W=480e-9 AD=76.8e-15 AS=76.8e-15 PD=1.26e-6 PS=1.26e-6 NRD=1.16667 NRS=1.16667 M=1
mi2__pm9 n215__vdd i2__net76 n10__i2__net77 n134__vdd g45p1svt L=45e-9 W=480e-9 AD=67.2e-15 AS=67.2e-15 PD=1.26e-6 PS=1.26e-6 NRD=1.16667 NRS=1.16667 M=1
mi2__pm11 n23__serial_out n4__i2__net77 n214__vdd n134__vdd g45p1svt L=45e-9 W=480e-9 AD=67.2e-15 AS=67.2e-15 PD=1.24e-6 PS=1.24e-6 NRD=1.16667 NRS=1.16667 M=1
mi2__pm13 i2__q n7__serial_out n213__vdd n134__vdd g45p1svt L=45e-9 W=480e-9 AD=67.2e-15 AS=67.2e-15 PD=1.24e-6 PS=1.24e-6 NRD=1.16667 NRS=1.16667 M=1
mi2__pm18 n9__i2__net79 shift n223__vdd n134__vdd g45p1svt L=45e-9 W=240e-9 AD=33.6e-15 AS=33.6e-15 PD=760e-9 PS=760e-9 NRD=1.16667 NRS=1.16667 M=1
mi2__pm16 n5__i2__net1 i2__net79 n4__net4 n134__vdd g45p1svt L=45e-9 W=240e-9 AD=38.4e-15 AS=38.4e-15 PD=780e-9 PS=780e-9 NRD=1.16667 NRS=1.16667 M=1
mi2__pm19 n3__r0_buff n20__shift n5__i2__net1 n134__vdd g45p1svt L=45e-9 W=240e-9 AD=33.6e-15 AS=33.6e-15 PD=780e-9 PS=780e-9 NRD=1.16667 NRS=1.16667 M=1
mi2__pm3 n6__i2__net73 i2__net1 n222__vdd n134__vdd g45p1svt L=45e-9 W=480e-9 AD=67.2e-15 AS=67.2e-15 PD=1.24e-6 PS=1.24e-6 NRD=1.16667 NRS=1.16667 M=1
mi2__pm0 n13__i2__net74 n17__ck_buff i2__net73 n134__vdd g45p1svt L=45e-9 W=120e-9 AD=16.8e-15 AS=16.8e-15 PD=520e-9 PS=520e-9 NRD=1.16667 NRS=1.16667 M=1
mi2__pm2 n221__vdd n3__i2__net75 n9__i2__net74 n134__vdd g45p1svt L=180e-9 W=120e-9 AD=16.8e-15 AS=16.8e-15 PD=520e-9 PS=520e-9 NRD=1.16667 NRS=1.16667 M=1
mi1__pm1_1__rcx n9__i1__net75 n6__i1__net74 n369__vdd n293__vdd g45p1svt L=45e-9 W=480e-9 AD=76.8e-15 AS=76.8e-15 PD=1.26e-6 PS=1.26e-6 NRD=1.16667 NRS=1.16667 M=1
mi1__pm1 n367__vdd n5__i1__net74 n9__i1__net75 n293__vdd g45p1svt L=45e-9 W=480e-9 AD=67.2e-15 AS=67.2e-15 PD=1.26e-6 PS=1.26e-6 NRD=1.16667 NRS=1.16667 M=1
mi1__pm8 n12__i1__net76 n28__ck_b n11__i1__net75 n293__vdd g45p1svt L=45e-9 W=120e-9 AD=16.8e-15 AS=16.8e-15 PD=520e-9 PS=520e-9 NRD=1.16667 NRS=1.16667 M=1
mi1__pm10 n365__vdd n2__i1__net77 n9__i1__net76 n293__vdd g45p1svt L=180e-9 W=120e-9 AD=16.8e-15 AS=16.8e-15 PD=520e-9 PS=520e-9 NRD=1.16667 NRS=1.16667 M=1
mi1__pm15 n15__i1__net76 n17__reset_b n363__vdd n293__vdd g45p1svt L=45e-9 W=120e-9 AD=16.8e-15 AS=16.8e-15 PD=520e-9 PS=520e-9 NRD=1.16667 NRS=1.16667 M=1
mi1__pm9_1__rcx n10__i1__net77 n6__i1__net76 n361__vdd n293__vdd g45p1svt L=45e-9 W=480e-9 AD=76.8e-15 AS=76.8e-15 PD=1.26e-6 PS=1.26e-6 NRD=1.16667 NRS=1.16667 M=1
mi1__pm9 n359__vdd n5__i1__net76 n10__i1__net77 n293__vdd g45p1svt L=45e-9 W=480e-9 AD=67.2e-15 AS=67.2e-15 PD=1.26e-6 PS=1.26e-6 NRD=1.16667 NRS=1.16667 M=1
mi1__pm11 n14__net4 n6__i1__net77 n357__vdd n293__vdd g45p1svt L=45e-9 W=480e-9 AD=67.2e-15 AS=67.2e-15 PD=1.24e-6 PS=1.24e-6 NRD=1.16667 NRS=1.16667 M=1
mi1__pm13 n3__i1__q n11__net4 n355__vdd n293__vdd g45p1svt L=45e-9 W=480e-9 AD=67.2e-15 AS=67.2e-15 PD=1.24e-6 PS=1.24e-6 NRD=1.16667 NRS=1.16667 M=1
mi1__pm18 n9__i1__net79 n8__shift n375__vdd n293__vdd g45p1svt L=45e-9 W=240e-9 AD=33.6e-15 AS=33.6e-15 PD=760e-9 PS=760e-9 NRD=1.16667 NRS=1.16667 M=1
mi1__pm16 n5__i1__net1 i1__net79 n4__net3 n293__vdd g45p1svt L=45e-9 W=240e-9 AD=38.4e-15 AS=38.4e-15 PD=780e-9 PS=780e-9 NRD=1.16667 NRS=1.16667 M=1
mi1__pm19 n3__r1_buff n22__shift n5__i1__net1 n293__vdd g45p1svt L=45e-9 W=240e-9 AD=33.6e-15 AS=33.6e-15 PD=780e-9 PS=780e-9 NRD=1.16667 NRS=1.16667 M=1
mi1__pm3 n4__i1__net73 n4__i1__net1 n373__vdd n293__vdd g45p1svt L=45e-9 W=480e-9 AD=67.2e-15 AS=67.2e-15 PD=1.24e-6 PS=1.24e-6 NRD=1.16667 NRS=1.16667 M=1
mi1__pm0 n12__i1__net74 n19__ck_buff n5__i1__net73 n293__vdd g45p1svt L=45e-9 W=120e-9 AD=16.8e-15 AS=16.8e-15 PD=520e-9 PS=520e-9 NRD=1.16667 NRS=1.16667 M=1
mi1__pm2 n371__vdd n2__i1__net75 n9__i1__net74 n293__vdd g45p1svt L=180e-9 W=120e-9 AD=16.8e-15 AS=16.8e-15 PD=520e-9 PS=520e-9 NRD=1.16667 NRS=1.16667 M=1
mi0__pm1_1__rcx n11__i0__net75 n7__i0__net74 n368__vdd n293__vdd g45p1svt L=45e-9 W=480e-9 AD=76.8e-15 AS=76.8e-15 PD=1.26e-6 PS=1.26e-6 NRD=1.16667 NRS=1.16667 M=1
mi0__pm1 n366__vdd i0__net74 n11__i0__net75 n293__vdd g45p1svt L=45e-9 W=480e-9 AD=67.2e-15 AS=67.2e-15 PD=1.26e-6 PS=1.26e-6 NRD=1.16667 NRS=1.16667 M=1
mi0__pm8 n13__i0__net76 n30__ck_b n6__i0__net75 n293__vdd g45p1svt L=45e-9 W=120e-9 AD=16.8e-15 AS=16.8e-15 PD=520e-9 PS=520e-9 NRD=1.16667 NRS=1.16667 M=1
mi0__pm10 n364__vdd n3__i0__net77 n9__i0__net76 n293__vdd g45p1svt L=180e-9 W=120e-9 AD=16.8e-15 AS=16.8e-15 PD=520e-9 PS=520e-9 NRD=1.16667 NRS=1.16667 M=1
mi0__pm15 n15__i0__net76 n19__reset_b n362__vdd n293__vdd g45p1svt L=45e-9 W=120e-9 AD=16.8e-15 AS=16.8e-15 PD=520e-9 PS=520e-9 NRD=1.16667 NRS=1.16667 M=1
mi0__pm9_1__rcx n10__i0__net77 n7__i0__net76 n360__vdd n293__vdd g45p1svt L=45e-9 W=480e-9 AD=76.8e-15 AS=76.8e-15 PD=1.26e-6 PS=1.26e-6 NRD=1.16667 NRS=1.16667 M=1
mi0__pm9 n358__vdd i0__net76 n10__i0__net77 n293__vdd g45p1svt L=45e-9 W=480e-9 AD=67.2e-15 AS=67.2e-15 PD=1.26e-6 PS=1.26e-6 NRD=1.16667 NRS=1.16667 M=1
mi0__pm11 n13__net3 n4__i0__net77 n356__vdd n293__vdd g45p1svt L=45e-9 W=480e-9 AD=67.2e-15 AS=67.2e-15 PD=1.24e-6 PS=1.24e-6 NRD=1.16667 NRS=1.16667 M=1
mi0__pm13 i0__q n6__net3 n354__vdd n293__vdd g45p1svt L=45e-9 W=480e-9 AD=67.2e-15 AS=67.2e-15 PD=1.24e-6 PS=1.24e-6 NRD=1.16667 NRS=1.16667 M=1
mi0__pm18 n9__i0__net79 n9__shift n374__vdd n293__vdd g45p1svt L=45e-9 W=240e-9 AD=33.6e-15 AS=33.6e-15 PD=760e-9 PS=760e-9 NRD=1.16667 NRS=1.16667 M=1
mi0__pm16 n5__i0__net1 i0__net79 n528__vss n293__vdd g45p1svt L=45e-9 W=240e-9 AD=38.4e-15 AS=38.4e-15 PD=780e-9 PS=780e-9 NRD=1.16667 NRS=1.16667 M=1
mi0__pm19 n3__r2_buff n24__shift n5__i0__net1 n293__vdd g45p1svt L=45e-9 W=240e-9 AD=33.6e-15 AS=33.6e-15 PD=780e-9 PS=780e-9 NRD=1.16667 NRS=1.16667 M=1
mi0__pm3 n6__i0__net73 i0__net1 n372__vdd n293__vdd g45p1svt L=45e-9 W=480e-9 AD=67.2e-15 AS=67.2e-15 PD=1.24e-6 PS=1.24e-6 NRD=1.16667 NRS=1.16667 M=1
mi0__pm0 n13__i0__net74 n21__ck_buff i0__net73 n293__vdd g45p1svt L=45e-9 W=120e-9 AD=16.8e-15 AS=16.8e-15 PD=520e-9 PS=520e-9 NRD=1.16667 NRS=1.16667 M=1
mi0__pm2 n370__vdd n3__i0__net75 n9__i0__net74 n293__vdd g45p1svt L=180e-9 W=120e-9 AD=16.8e-15 AS=16.8e-15 PD=520e-9 PS=520e-9 NRD=1.16667 NRS=1.16667 M=1
mi14__pm2_5__rcx n249__vdd n22__i14__net7 n88__i14__net9 n134__vdd g45p1svt L=45e-9 W=480e-9 AD=76.8e-15 AS=76.8e-15 PD=1.28e-6 PS=1.28e-6 NRD=1.16667 NRS=1.16667 M=1
mi14__pm2_4__rcx n91__i14__net9 n20__i14__net7 n249__vdd n134__vdd g45p1svt L=45e-9 W=480e-9 AD=76.8e-15 AS=76.8e-15 PD=1.28e-6 PS=1.28e-6 NRD=1.16667 NRS=1.16667 M=1
mi14__pm2_3__rcx n247__vdd n18__i14__net7 n91__i14__net9 n134__vdd g45p1svt L=45e-9 W=480e-9 AD=76.8e-15 AS=76.8e-15 PD=1.28e-6 PS=1.28e-6 NRD=1.16667 NRS=1.16667 M=1
mi14__pm2_2__rcx n94__i14__net9 n16__i14__net7 n247__vdd n134__vdd g45p1svt L=45e-9 W=480e-9 AD=76.8e-15 AS=76.8e-15 PD=1.28e-6 PS=1.28e-6 NRD=1.16667 NRS=1.16667 M=1
mi14__pm2_1__rcx n245__vdd n15__i14__net7 n94__i14__net9 n134__vdd g45p1svt L=45e-9 W=480e-9 AD=67.2e-15 AS=67.2e-15 PD=1.26e-6 PS=1.26e-6 NRD=1.16667 NRS=1.16667 M=1
mi14__pm2 n88__i14__net9 n14__i14__net7 n251__vdd n134__vdd g45p1svt L=45e-9 W=480e-9 AD=76.8e-15 AS=76.8e-15 PD=1.26e-6 PS=1.26e-6 NRD=1.16667 NRS=1.16667 M=1
mi14__pm8_5__rcx n264__vdd n43__reset n51__i14__net4 n134__vdd g45p1svt L=45e-9 W=480e-9 AD=76.8e-15 AS=76.8e-15 PD=1.28e-6 PS=1.28e-6 NRD=1.16667 NRS=1.16667 M=1
mi14__pm8_4__rcx n54__i14__net4 n41__reset n264__vdd n134__vdd g45p1svt L=45e-9 W=480e-9 AD=76.8e-15 AS=76.8e-15 PD=1.28e-6 PS=1.28e-6 NRD=1.16667 NRS=1.16667 M=1
mi14__pm8_3__rcx n259__vdd n39__reset n54__i14__net4 n134__vdd g45p1svt L=45e-9 W=480e-9 AD=76.8e-15 AS=76.8e-15 PD=1.28e-6 PS=1.28e-6 NRD=1.16667 NRS=1.16667 M=1
mi14__pm8_2__rcx n57__i14__net4 n37__reset n259__vdd n134__vdd g45p1svt L=45e-9 W=480e-9 AD=76.8e-15 AS=76.8e-15 PD=1.28e-6 PS=1.28e-6 NRD=1.16667 NRS=1.16667 M=1
mi14__pm8_1__rcx n258__vdd n36__reset n57__i14__net4 n134__vdd g45p1svt L=45e-9 W=480e-9 AD=67.2e-15 AS=67.2e-15 PD=1.26e-6 PS=1.26e-6 NRD=1.16667 NRS=1.16667 M=1
mi14__pm8 n51__i14__net4 n35__reset n265__vdd n134__vdd g45p1svt L=45e-9 W=480e-9 AD=76.8e-15 AS=76.8e-15 PD=1.26e-6 PS=1.26e-6 NRD=1.16667 NRS=1.16667 M=1
mi14__pm3_5__rcx n248__vdd n23__i14__net11 n97__i14__net10 n134__vdd g45p1svt L=45e-9 W=480e-9 AD=76.8e-15 AS=76.8e-15 PD=1.28e-6 PS=1.28e-6 NRD=1.16667 NRS=1.16667 M=1
mi14__pm3_4__rcx n100__i14__net10 n21__i14__net11 n248__vdd n134__vdd g45p1svt L=45e-9 W=480e-9 AD=76.8e-15 AS=76.8e-15 PD=1.28e-6 PS=1.28e-6 NRD=1.16667 NRS=1.16667 M=1
mi14__pm3_3__rcx n246__vdd n19__i14__net11 n100__i14__net10 n134__vdd g45p1svt L=45e-9 W=480e-9 AD=76.8e-15 AS=76.8e-15 PD=1.28e-6 PS=1.28e-6 NRD=1.16667 NRS=1.16667 M=1
mi14__pm3_2__rcx n103__i14__net10 n17__i14__net11 n246__vdd n134__vdd g45p1svt L=45e-9 W=480e-9 AD=76.8e-15 AS=76.8e-15 PD=1.28e-6 PS=1.28e-6 NRD=1.16667 NRS=1.16667 M=1
mi14__pm3_1__rcx n244__vdd n5__i14__net11 n103__i14__net10 n134__vdd g45p1svt L=45e-9 W=480e-9 AD=67.2e-15 AS=67.2e-15 PD=1.26e-6 PS=1.26e-6 NRD=1.16667 NRS=1.16667 M=1
mi14__pm3 n97__i14__net10 n24__i14__net11 n250__vdd n134__vdd g45p1svt L=45e-9 W=480e-9 AD=76.8e-15 AS=76.8e-15 PD=1.26e-6 PS=1.26e-6 NRD=1.16667 NRS=1.16667 M=1
mi14__pm7_5__rcx n256__vdd n47__i14__net4 n57__i14__net3 n134__vdd g45p1svt L=45e-9 W=480e-9 AD=76.8e-15 AS=76.8e-15 PD=1.28e-6 PS=1.28e-6 NRD=1.16667 NRS=1.16667 M=1
mi14__pm7_4__rcx n60__i14__net3 n45__i14__net4 n256__vdd n134__vdd g45p1svt L=45e-9 W=480e-9 AD=76.8e-15 AS=76.8e-15 PD=1.28e-6 PS=1.28e-6 NRD=1.16667 NRS=1.16667 M=1
mi14__pm7_3__rcx n254__vdd n43__i14__net4 n60__i14__net3 n134__vdd g45p1svt L=45e-9 W=480e-9 AD=76.8e-15 AS=76.8e-15 PD=1.28e-6 PS=1.28e-6 NRD=1.16667 NRS=1.16667 M=1
mi14__pm7_2__rcx n70__i14__net3 n41__i14__net4 n254__vdd n134__vdd g45p1svt L=45e-9 W=480e-9 AD=76.8e-15 AS=76.8e-15 PD=1.28e-6 PS=1.28e-6 NRD=1.16667 NRS=1.16667 M=1
mi14__pm7_1__rcx n252__vdd n29__i14__net4 n70__i14__net3 n134__vdd g45p1svt L=45e-9 W=480e-9 AD=67.2e-15 AS=67.2e-15 PD=1.26e-6 PS=1.26e-6 NRD=1.16667 NRS=1.16667 M=1
mi14__pm7 n57__i14__net3 n48__i14__net4 n257__vdd n134__vdd g45p1svt L=45e-9 W=480e-9 AD=76.8e-15 AS=76.8e-15 PD=1.26e-6 PS=1.26e-6 NRD=1.16667 NRS=1.16667 M=1
mi14__i17__i2__pm0 n12__i14__i17__i2__net1 n5__ck n7__i14__i17__net1 n134__vdd g45p1svt L=45e-9 W=120e-9 AD=16.8e-15 AS=16.8e-15 PD=520e-9 PS=520e-9 NRD=1.16667 NRS=1.16667 M=1
mi14__i17__i2__pm2 n289__vdd n2__i14__i17__i2__net2 n9__i14__i17__i2__net1 n134__vdd g45p1svt L=180e-9 W=120e-9 AD=16.8e-15 AS=16.8e-15 PD=520e-9 PS=520e-9 NRD=1.16667 NRS=1.16667 M=1
mi14__i17__i2__pm1_1__rcx n9__i14__i17__i2__net2 n6__i14__i17__i2__net1 n287__vdd n134__vdd g45p1svt L=45e-9 W=480e-9 AD=76.8e-15 AS=76.8e-15 PD=1.26e-6 PS=1.26e-6 NRD=1.16667 NRS=1.16667 M=1
mi14__i17__i2__pm1 n285__vdd n5__i14__i17__i2__net1 n9__i14__i17__i2__net2 n134__vdd g45p1svt L=45e-9 W=480e-9 AD=67.2e-15 AS=67.2e-15 PD=1.26e-6 PS=1.26e-6 NRD=1.16667 NRS=1.16667 M=1
mi14__i17__i2__pm8 n12__i14__i17__i2__net5 n4__i14__i17__net3 n11__i14__i17__i2__net2 n134__vdd g45p1svt L=45e-9 W=120e-9 AD=16.8e-15 AS=16.8e-15 PD=520e-9 PS=520e-9 NRD=1.16667 NRS=1.16667 M=1
mi14__i17__i2__pm10 n283__vdd n2__i14__i17__i2__net4 n9__i14__i17__i2__net5 n134__vdd g45p1svt L=180e-9 W=120e-9 AD=16.8e-15 AS=16.8e-15 PD=520e-9 PS=520e-9 NRD=1.16667 NRS=1.16667 M=1
mi14__i17__i2__pm15 n15__i14__i17__i2__net5 i14__i17__net6 n281__vdd n134__vdd g45p1svt L=45e-9 W=120e-9 AD=16.8e-15 AS=16.8e-15 PD=520e-9 PS=520e-9 NRD=1.16667 NRS=1.16667 M=1
mi14__i17__i2__pm9_1__rcx n10__i14__i17__i2__net4 n6__i14__i17__i2__net5 n279__vdd n134__vdd g45p1svt L=45e-9 W=480e-9 AD=76.8e-15 AS=76.8e-15 PD=1.26e-6 PS=1.26e-6 NRD=1.16667 NRS=1.16667 M=1
mi14__i17__i2__pm9 n277__vdd n5__i14__i17__i2__net5 n10__i14__i17__i2__net4 n134__vdd g45p1svt L=45e-9 W=480e-9 AD=67.2e-15 AS=67.2e-15 PD=1.26e-6 PS=1.26e-6 NRD=1.16667 NRS=1.16667 M=1
mi14__i17__i2__pm11 n28__i14__i17__net1 n6__i14__i17__i2__net4 n275__vdd n134__vdd g45p1svt L=45e-9 W=480e-9 AD=67.2e-15 AS=67.2e-15 PD=1.24e-6 PS=1.24e-6 NRD=1.16667 NRS=1.16667 M=1
mi14__i17__i2__pm13 n19__i14__i17__net7 n17__i14__i17__net1 n273__vdd n134__vdd g45p1svt L=45e-9 W=480e-9 AD=67.2e-15 AS=67.2e-15 PD=1.24e-6 PS=1.24e-6 NRD=1.16667 NRS=1.16667 M=1
mi14__i17__i3__pm0 n13__i14__i17__i3__net1 n2__i14__i17__net7 i14__i17__net8 n134__vdd g45p1svt L=45e-9 W=120e-9 AD=16.8e-15 AS=16.8e-15 PD=520e-9 PS=520e-9 NRD=1.16667 NRS=1.16667 M=1
mi14__i17__i3__pm2 n288__vdd n3__i14__i17__i3__net2 n9__i14__i17__i3__net1 n134__vdd g45p1svt L=180e-9 W=120e-9 AD=16.8e-15 AS=16.8e-15 PD=520e-9 PS=520e-9 NRD=1.16667 NRS=1.16667 M=1
mi14__i17__i3__pm1_1__rcx n11__i14__i17__i3__net2 n7__i14__i17__i3__net1 n286__vdd n134__vdd g45p1svt L=45e-9 W=480e-9 AD=76.8e-15 AS=76.8e-15 PD=1.26e-6 PS=1.26e-6 NRD=1.16667 NRS=1.16667 M=1
mi14__i17__i3__pm1 n284__vdd i14__i17__i3__net1 n11__i14__i17__i3__net2 n134__vdd g45p1svt L=45e-9 W=480e-9 AD=67.2e-15 AS=67.2e-15 PD=1.26e-6 PS=1.26e-6 NRD=1.16667 NRS=1.16667 M=1
mi14__i17__i3__pm8 n13__i14__i17__i3__net5 n4__i14__i17__net1 n6__i14__i17__i3__net2 n134__vdd g45p1svt L=45e-9 W=120e-9 AD=16.8e-15 AS=16.8e-15 PD=520e-9 PS=520e-9 NRD=1.16667 NRS=1.16667 M=1
mi14__i17__i3__pm10 n282__vdd n3__i14__i17__i3__net4 n9__i14__i17__i3__net5 n134__vdd g45p1svt L=180e-9 W=120e-9 AD=16.8e-15 AS=16.8e-15 PD=520e-9 PS=520e-9 NRD=1.16667 NRS=1.16667 M=1
mi14__i17__i3__pm15 n15__i14__i17__i3__net5 n3__i14__i17__net6 n280__vdd n134__vdd g45p1svt L=45e-9 W=120e-9 AD=16.8e-15 AS=16.8e-15 PD=520e-9 PS=520e-9 NRD=1.16667 NRS=1.16667 M=1
mi14__i17__i3__pm9_1__rcx n10__i14__i17__i3__net4 n7__i14__i17__i3__net5 n278__vdd n134__vdd g45p1svt L=45e-9 W=480e-9 AD=76.8e-15 AS=76.8e-15 PD=1.26e-6 PS=1.26e-6 NRD=1.16667 NRS=1.16667 M=1
mi14__i17__i3__pm9 n276__vdd i14__i17__i3__net5 n10__i14__i17__i3__net4 n134__vdd g45p1svt L=45e-9 W=480e-9 AD=67.2e-15 AS=67.2e-15 PD=1.26e-6 PS=1.26e-6 NRD=1.16667 NRS=1.16667 M=1
mi14__i17__i3__pm11 n22__i14__i17__net8 n4__i14__i17__i3__net4 n274__vdd n134__vdd g45p1svt L=45e-9 W=480e-9 AD=67.2e-15 AS=67.2e-15 PD=1.24e-6 PS=1.24e-6 NRD=1.16667 NRS=1.16667 M=1
mi14__i17__i3__pm13 n10__i14__i17__net11 n6__i14__i17__net8 n272__vdd n134__vdd g45p1svt L=45e-9 W=480e-9 AD=67.2e-15 AS=67.2e-15 PD=1.24e-6 PS=1.24e-6 NRD=1.16667 NRS=1.16667 M=1
mi14__i17__i4__pm3 n8__i14__i17__net9 n10__i14__i17__net8 n853__vss n134__vdd g45p1svt L=45e-9 W=240e-9 AD=38.4e-15 AS=38.4e-15 PD=780e-9 PS=780e-9 NRD=1.16667 NRS=1.16667 M=1
mi14__i17__i4__pm2 n268__vdd n2__i14__i17__net11 n8__i14__i17__net9 n134__vdd g45p1svt L=45e-9 W=240e-9 AD=33.6e-15 AS=33.6e-15 PD=780e-9 PS=780e-9 NRD=1.16667 NRS=1.16667 M=1
mi14__i17__i4__pm6 n11__i14__i17__net10 n5__i14__i17__net9 n266__vdd n134__vdd g45p1svt L=45e-9 W=480e-9 AD=67.2e-15 AS=67.2e-15 PD=1.24e-6 PS=1.24e-6 NRD=1.16667 NRS=1.16667 M=1
mi14__i17__i4__pm5 n263__vdd n5__i14__i17__net10 n18__i14__i17__net9 n134__vdd g45p1svt L=45e-9 W=480e-9 AD=67.2e-15 AS=67.2e-15 PD=1.24e-6 PS=1.24e-6 NRD=1.16667 NRS=1.16667 M=1
mi14__i17__i4__pm0 n18__i14__i17__net10 n15__i14__i17__net8 n260__vdd n134__vdd g45p1svt L=45e-9 W=240e-9 AD=38.4e-15 AS=38.4e-15 PD=780e-9 PS=780e-9 NRD=1.16667 NRS=1.16667 M=1
mi14__i17__i4__pm1 n837__vss n6__i14__i17__net11 n18__i14__i17__net10 n134__vdd g45p1svt L=45e-9 W=240e-9 AD=33.6e-15 AS=33.6e-15 PD=780e-9 PS=780e-9 NRD=1.16667 NRS=1.16667 M=1
mi14__i17__pm17 n25__i14__net7 n4__i14__i17__net9 n267__vdd n134__vdd g45p1svt L=45e-9 W=480e-9 AD=67.2e-15 AS=67.2e-15 PD=1.24e-6 PS=1.24e-6 NRD=1.16667 NRS=1.16667 M=1
mi14__i17__pm16 n26__i14__net11 n4__i14__i17__net10 n271__vdd n134__vdd g45p1svt L=45e-9 W=480e-9 AD=67.2e-15 AS=67.2e-15 PD=1.24e-6 PS=1.24e-6 NRD=1.16667 NRS=1.16667 M=1
mi14__i17__pm1 n5__i14__i17__net6 n1__reset n210__vdd n134__vdd g45p1svt L=45e-9 W=240e-9 AD=33.6e-15 AS=33.6e-15 PD=760e-9 PS=760e-9 NRD=1.16667 NRS=1.16667 M=1
mi14__i17__pm0 n7__i14__i17__net3 n3__ck n290__vdd n134__vdd g45p1svt L=45e-9 W=240e-9 AD=33.6e-15 AS=33.6e-15 PD=760e-9 PS=760e-9 NRD=1.16667 NRS=1.16667 M=1
mi14__i11__pm0 n12__i14__i11__net1 n30__i14__net10 n3__y3 n293__vdd g45p1svt L=45e-9 W=120e-9 AD=16.8e-15 AS=16.8e-15 PD=520e-9 PS=520e-9 NRD=1.16667 NRS=1.16667 M=1
mi14__i11__pm2 n401__vdd n2__i14__i11__net2 n9__i14__i11__net1 n293__vdd g45p1svt L=180e-9 W=120e-9 AD=16.8e-15 AS=16.8e-15 PD=520e-9 PS=520e-9 NRD=1.16667 NRS=1.16667 M=1
mi14__i11__pm1_1__rcx n9__i14__i11__net2 n6__i14__i11__net1 n399__vdd n293__vdd g45p1svt L=45e-9 W=480e-9 AD=76.8e-15 AS=76.8e-15 PD=1.26e-6 PS=1.26e-6 NRD=1.16667 NRS=1.16667 M=1
mi14__i11__pm1 n397__vdd n5__i14__i11__net1 n9__i14__i11__net2 n293__vdd g45p1svt L=45e-9 W=480e-9 AD=67.2e-15 AS=67.2e-15 PD=1.26e-6 PS=1.26e-6 NRD=1.16667 NRS=1.16667 M=1
mi14__i11__pm8 n12__i14__i11__net5 n50__i14__net9 n11__i14__i11__net2 n293__vdd g45p1svt L=45e-9 W=120e-9 AD=16.8e-15 AS=16.8e-15 PD=520e-9 PS=520e-9 NRD=1.16667 NRS=1.16667 M=1
mi14__i11__pm10 n395__vdd n2__i14__i11__net4 n9__i14__i11__net5 n293__vdd g45p1svt L=180e-9 W=120e-9 AD=16.8e-15 AS=16.8e-15 PD=520e-9 PS=520e-9 NRD=1.16667 NRS=1.16667 M=1
mi14__i11__pm15 n15__i14__i11__net5 n21__i14__net4 n393__vdd n293__vdd g45p1svt L=45e-9 W=120e-9 AD=16.8e-15 AS=16.8e-15 PD=520e-9 PS=520e-9 NRD=1.16667 NRS=1.16667 M=1
mi14__i11__pm9_1__rcx n11__i14__i11__net4 n6__i14__i11__net5 n391__vdd n293__vdd g45p1svt L=45e-9 W=480e-9 AD=76.8e-15 AS=76.8e-15 PD=1.26e-6 PS=1.26e-6 NRD=1.16667 NRS=1.16667 M=1
mi14__i11__pm9 n389__vdd n5__i14__i11__net5 n11__i14__i11__net4 n293__vdd g45p1svt L=45e-9 W=480e-9 AD=67.2e-15 AS=67.2e-15 PD=1.26e-6 PS=1.26e-6 NRD=1.16667 NRS=1.16667 M=1
mi14__i11__pm11 n9__i14__x_out_b_1 n6__i14__i11__net4 n387__vdd n293__vdd g45p1svt L=45e-9 W=480e-9 AD=67.2e-15 AS=67.2e-15 PD=1.24e-6 PS=1.24e-6 NRD=1.16667 NRS=1.16667 M=1
mi14__i11__pm13 n9__y_out_3 n4__i14__x_out_b_1 n385__vdd n293__vdd g45p1svt L=45e-9 W=480e-9 AD=67.2e-15 AS=67.2e-15 PD=1.24e-6 PS=1.24e-6 NRD=1.16667 NRS=1.16667 M=1
mi14__i13__pm0 n12__i14__i13__net1 n2__i14__net10 n3__x3 n293__vdd g45p1svt L=45e-9 W=120e-9 AD=16.8e-15 AS=16.8e-15 PD=520e-9 PS=520e-9 NRD=1.16667 NRS=1.16667 M=1
mi14__i13__pm2 n418__vdd n2__i14__i13__net2 n9__i14__i13__net1 n293__vdd g45p1svt L=180e-9 W=120e-9 AD=16.8e-15 AS=16.8e-15 PD=520e-9 PS=520e-9 NRD=1.16667 NRS=1.16667 M=1
mi14__i13__pm1_1__rcx n9__i14__i13__net2 n6__i14__i13__net1 n417__vdd n293__vdd g45p1svt L=45e-9 W=480e-9 AD=76.8e-15 AS=76.8e-15 PD=1.26e-6 PS=1.26e-6 NRD=1.16667 NRS=1.16667 M=1
mi14__i13__pm1 n415__vdd n5__i14__i13__net1 n9__i14__i13__net2 n293__vdd g45p1svt L=45e-9 W=480e-9 AD=67.2e-15 AS=67.2e-15 PD=1.26e-6 PS=1.26e-6 NRD=1.16667 NRS=1.16667 M=1
mi14__i13__pm8 n12__i14__i13__net5 n10__i14__net9 n11__i14__i13__net2 n293__vdd g45p1svt L=45e-9 W=120e-9 AD=16.8e-15 AS=16.8e-15 PD=520e-9 PS=520e-9 NRD=1.16667 NRS=1.16667 M=1
mi14__i13__pm10 n413__vdd n2__i14__i13__net4 n9__i14__i13__net5 n293__vdd g45p1svt L=180e-9 W=120e-9 AD=16.8e-15 AS=16.8e-15 PD=520e-9 PS=520e-9 NRD=1.16667 NRS=1.16667 M=1
mi14__i13__pm15 n15__i14__i13__net5 i14__net4 n411__vdd n293__vdd g45p1svt L=45e-9 W=120e-9 AD=16.8e-15 AS=16.8e-15 PD=520e-9 PS=520e-9 NRD=1.16667 NRS=1.16667 M=1
mi14__i13__pm9_1__rcx n10__i14__i13__net4 n6__i14__i13__net5 n409__vdd n293__vdd g45p1svt L=45e-9 W=480e-9 AD=76.8e-15 AS=76.8e-15 PD=1.26e-6 PS=1.26e-6 NRD=1.16667 NRS=1.16667 M=1
mi14__i13__pm9 n407__vdd n5__i14__i13__net5 n10__i14__i13__net4 n293__vdd g45p1svt L=45e-9 W=480e-9 AD=67.2e-15 AS=67.2e-15 PD=1.26e-6 PS=1.26e-6 NRD=1.16667 NRS=1.16667 M=1
mi14__i13__pm11 n9__i14__y_out_b_3 n6__i14__i13__net4 n405__vdd n293__vdd g45p1svt L=45e-9 W=480e-9 AD=67.2e-15 AS=67.2e-15 PD=1.24e-6 PS=1.24e-6 NRD=1.16667 NRS=1.16667 M=1
mi14__i13__pm13 n3__x_out_3 n4__i14__y_out_b_3 n403__vdd n293__vdd g45p1svt L=45e-9 W=480e-9 AD=67.2e-15 AS=67.2e-15 PD=1.24e-6 PS=1.24e-6 NRD=1.16667 NRS=1.16667 M=1
mi14__i15__pm0 n12__i14__i15__net1 n34__i14__net10 n3__y1 n32__vdd g45p1svt L=45e-9 W=120e-9 AD=16.8e-15 AS=16.8e-15 PD=520e-9 PS=520e-9 NRD=1.16667 NRS=1.16667 M=1
mi14__i15__pm2 n106__vdd n2__i14__i15__net2 n9__i14__i15__net1 n32__vdd g45p1svt L=180e-9 W=120e-9 AD=16.8e-15 AS=16.8e-15 PD=520e-9 PS=520e-9 NRD=1.16667 NRS=1.16667 M=1
mi14__i15__pm1_1__rcx n9__i14__i15__net2 n6__i14__i15__net1 n104__vdd n32__vdd g45p1svt L=45e-9 W=480e-9 AD=76.8e-15 AS=76.8e-15 PD=1.26e-6 PS=1.26e-6 NRD=1.16667 NRS=1.16667 M=1
mi14__i15__pm1 n102__vdd n5__i14__i15__net1 n9__i14__i15__net2 n32__vdd g45p1svt L=45e-9 W=480e-9 AD=67.2e-15 AS=67.2e-15 PD=1.26e-6 PS=1.26e-6 NRD=1.16667 NRS=1.16667 M=1
mi14__i15__pm8 n12__i14__i15__net5 n54__i14__net9 n11__i14__i15__net2 n32__vdd g45p1svt L=45e-9 W=120e-9 AD=16.8e-15 AS=16.8e-15 PD=520e-9 PS=520e-9 NRD=1.16667 NRS=1.16667 M=1
mi14__i15__pm10 n100__vdd n2__i14__i15__net4 n9__i14__i15__net5 n32__vdd g45p1svt L=180e-9 W=120e-9 AD=16.8e-15 AS=16.8e-15 PD=520e-9 PS=520e-9 NRD=1.16667 NRS=1.16667 M=1
mi14__i15__pm15 n15__i14__i15__net5 n25__i14__net4 n98__vdd n32__vdd g45p1svt L=45e-9 W=120e-9 AD=16.8e-15 AS=16.8e-15 PD=520e-9 PS=520e-9 NRD=1.16667 NRS=1.16667 M=1
mi14__i15__pm9_1__rcx n11__i14__i15__net4 n6__i14__i15__net5 n96__vdd n32__vdd g45p1svt L=45e-9 W=480e-9 AD=76.8e-15 AS=76.8e-15 PD=1.26e-6 PS=1.26e-6 NRD=1.16667 NRS=1.16667 M=1
mi14__i15__pm9 n94__vdd n5__i14__i15__net5 n11__i14__i15__net4 n32__vdd g45p1svt L=45e-9 W=480e-9 AD=67.2e-15 AS=67.2e-15 PD=1.26e-6 PS=1.26e-6 NRD=1.16667 NRS=1.16667 M=1
mi14__i15__pm11 n9__i14__y_out_b_1 n6__i14__i15__net4 n92__vdd n32__vdd g45p1svt L=45e-9 W=480e-9 AD=67.2e-15 AS=67.2e-15 PD=1.24e-6 PS=1.24e-6 NRD=1.16667 NRS=1.16667 M=1
mi14__i15__pm13 n9__y_out_1 n4__i14__y_out_b_1 n90__vdd n32__vdd g45p1svt L=45e-9 W=480e-9 AD=67.2e-15 AS=67.2e-15 PD=1.24e-6 PS=1.24e-6 NRD=1.16667 NRS=1.16667 M=1
mi14__i10__pm0 n12__i14__i10__net1 n6__i14__net10 n3__x1 n32__vdd g45p1svt L=45e-9 W=120e-9 AD=16.8e-15 AS=16.8e-15 PD=520e-9 PS=520e-9 NRD=1.16667 NRS=1.16667 M=1
mi14__i10__pm2 n129__vdd n2__i14__i10__net2 n9__i14__i10__net1 n32__vdd g45p1svt L=180e-9 W=120e-9 AD=16.8e-15 AS=16.8e-15 PD=520e-9 PS=520e-9 NRD=1.16667 NRS=1.16667 M=1
mi14__i10__pm1_1__rcx n9__i14__i10__net2 n6__i14__i10__net1 n127__vdd n32__vdd g45p1svt L=45e-9 W=480e-9 AD=76.8e-15 AS=76.8e-15 PD=1.26e-6 PS=1.26e-6 NRD=1.16667 NRS=1.16667 M=1
mi14__i10__pm1 n123__vdd n5__i14__i10__net1 n9__i14__i10__net2 n32__vdd g45p1svt L=45e-9 W=480e-9 AD=67.2e-15 AS=67.2e-15 PD=1.26e-6 PS=1.26e-6 NRD=1.16667 NRS=1.16667 M=1
mi14__i10__pm8 n12__i14__i10__net5 n14__i14__net9 n11__i14__i10__net2 n32__vdd g45p1svt L=45e-9 W=120e-9 AD=16.8e-15 AS=16.8e-15 PD=520e-9 PS=520e-9 NRD=1.16667 NRS=1.16667 M=1
mi14__i10__pm10 n120__vdd n2__i14__i10__net4 n9__i14__i10__net5 n32__vdd g45p1svt L=180e-9 W=120e-9 AD=16.8e-15 AS=16.8e-15 PD=520e-9 PS=520e-9 NRD=1.16667 NRS=1.16667 M=1
mi14__i10__pm15 n15__i14__i10__net5 n5__i14__net4 n116__vdd n32__vdd g45p1svt L=45e-9 W=120e-9 AD=16.8e-15 AS=16.8e-15 PD=520e-9 PS=520e-9 NRD=1.16667 NRS=1.16667 M=1
mi14__i10__pm9_1__rcx n10__i14__i10__net4 n6__i14__i10__net5 n114__vdd n32__vdd g45p1svt L=45e-9 W=480e-9 AD=76.8e-15 AS=76.8e-15 PD=1.26e-6 PS=1.26e-6 NRD=1.16667 NRS=1.16667 M=1
mi14__i10__pm9 n112__vdd n5__i14__i10__net5 n10__i14__i10__net4 n32__vdd g45p1svt L=45e-9 W=480e-9 AD=67.2e-15 AS=67.2e-15 PD=1.26e-6 PS=1.26e-6 NRD=1.16667 NRS=1.16667 M=1
mi14__i10__pm11 n9__i14__x_out_b_2 n6__i14__i10__net4 n110__vdd n32__vdd g45p1svt L=45e-9 W=480e-9 AD=67.2e-15 AS=67.2e-15 PD=1.24e-6 PS=1.24e-6 NRD=1.16667 NRS=1.16667 M=1
mi14__i10__pm13 n3__x_out_1 n4__i14__x_out_b_2 n108__vdd n32__vdd g45p1svt L=45e-9 W=480e-9 AD=67.2e-15 AS=67.2e-15 PD=1.24e-6 PS=1.24e-6 NRD=1.16667 NRS=1.16667 M=1
mi14__i14__pm0 n13__i14__i14__net1 n32__i14__net10 n1__y2 n293__vdd g45p1svt L=45e-9 W=120e-9 AD=16.8e-15 AS=16.8e-15 PD=520e-9 PS=520e-9 NRD=1.16667 NRS=1.16667 M=1
mi14__i14__pm2 n400__vdd n3__i14__i14__net2 n9__i14__i14__net1 n293__vdd g45p1svt L=180e-9 W=120e-9 AD=16.8e-15 AS=16.8e-15 PD=520e-9 PS=520e-9 NRD=1.16667 NRS=1.16667 M=1
mi14__i14__pm1_1__rcx n11__i14__i14__net2 n7__i14__i14__net1 n398__vdd n293__vdd g45p1svt L=45e-9 W=480e-9 AD=76.8e-15 AS=76.8e-15 PD=1.26e-6 PS=1.26e-6 NRD=1.16667 NRS=1.16667 M=1
mi14__i14__pm1 n396__vdd i14__i14__net1 n11__i14__i14__net2 n293__vdd g45p1svt L=45e-9 W=480e-9 AD=67.2e-15 AS=67.2e-15 PD=1.26e-6 PS=1.26e-6 NRD=1.16667 NRS=1.16667 M=1
mi14__i14__pm8 n13__i14__i14__net5 n52__i14__net9 n6__i14__i14__net2 n293__vdd g45p1svt L=45e-9 W=120e-9 AD=16.8e-15 AS=16.8e-15 PD=520e-9 PS=520e-9 NRD=1.16667 NRS=1.16667 M=1
mi14__i14__pm10 n394__vdd n3__i14__i14__net4 n9__i14__i14__net5 n293__vdd g45p1svt L=180e-9 W=120e-9 AD=16.8e-15 AS=16.8e-15 PD=520e-9 PS=520e-9 NRD=1.16667 NRS=1.16667 M=1
mi14__i14__pm15 n15__i14__i14__net5 n23__i14__net4 n392__vdd n293__vdd g45p1svt L=45e-9 W=120e-9 AD=16.8e-15 AS=16.8e-15 PD=520e-9 PS=520e-9 NRD=1.16667 NRS=1.16667 M=1
mi14__i14__pm9_1__rcx n11__i14__i14__net4 n7__i14__i14__net5 n390__vdd n293__vdd g45p1svt L=45e-9 W=480e-9 AD=76.8e-15 AS=76.8e-15 PD=1.26e-6 PS=1.26e-6 NRD=1.16667 NRS=1.16667 M=1
mi14__i14__pm9 n388__vdd i14__i14__net5 n11__i14__i14__net4 n293__vdd g45p1svt L=45e-9 W=480e-9 AD=67.2e-15 AS=67.2e-15 PD=1.26e-6 PS=1.26e-6 NRD=1.16667 NRS=1.16667 M=1
mi14__i14__pm11 n10__i14__y_out_b_2 n4__i14__i14__net4 n386__vdd n293__vdd g45p1svt L=45e-9 W=480e-9 AD=67.2e-15 AS=67.2e-15 PD=1.24e-6 PS=1.24e-6 NRD=1.16667 NRS=1.16667 M=1
mi14__i14__pm13 n7__y_out_2 i14__y_out_b_2 n384__vdd n293__vdd g45p1svt L=45e-9 W=480e-9 AD=67.2e-15 AS=67.2e-15 PD=1.24e-6 PS=1.24e-6 NRD=1.16667 NRS=1.16667 M=1
mi14__i16__pm0 n13__i14__i16__net1 n4__i14__net10 n1__x2 n293__vdd g45p1svt L=45e-9 W=120e-9 AD=16.8e-15 AS=16.8e-15 PD=520e-9 PS=520e-9 NRD=1.16667 NRS=1.16667 M=1
mi14__i16__pm2 n348__vdd n3__i14__i16__net2 n9__i14__i16__net1 n293__vdd g45p1svt L=180e-9 W=120e-9 AD=16.8e-15 AS=16.8e-15 PD=520e-9 PS=520e-9 NRD=1.16667 NRS=1.16667 M=1
mi14__i16__pm1_1__rcx n11__i14__i16__net2 n7__i14__i16__net1 n416__vdd n293__vdd g45p1svt L=45e-9 W=480e-9 AD=76.8e-15 AS=76.8e-15 PD=1.26e-6 PS=1.26e-6 NRD=1.16667 NRS=1.16667 M=1
mi14__i16__pm1 n414__vdd i14__i16__net1 n11__i14__i16__net2 n293__vdd g45p1svt L=45e-9 W=480e-9 AD=67.2e-15 AS=67.2e-15 PD=1.26e-6 PS=1.26e-6 NRD=1.16667 NRS=1.16667 M=1
mi14__i16__pm8 n13__i14__i16__net5 n12__i14__net9 n6__i14__i16__net2 n293__vdd g45p1svt L=45e-9 W=120e-9 AD=16.8e-15 AS=16.8e-15 PD=520e-9 PS=520e-9 NRD=1.16667 NRS=1.16667 M=1
mi14__i16__pm10 n412__vdd n3__i14__i16__net4 n9__i14__i16__net5 n293__vdd g45p1svt L=180e-9 W=120e-9 AD=16.8e-15 AS=16.8e-15 PD=520e-9 PS=520e-9 NRD=1.16667 NRS=1.16667 M=1
mi14__i16__pm15 n15__i14__i16__net5 n3__i14__net4 n410__vdd n293__vdd g45p1svt L=45e-9 W=120e-9 AD=16.8e-15 AS=16.8e-15 PD=520e-9 PS=520e-9 NRD=1.16667 NRS=1.16667 M=1
mi14__i16__pm9_1__rcx n10__i14__i16__net4 n7__i14__i16__net5 n408__vdd n293__vdd g45p1svt L=45e-9 W=480e-9 AD=76.8e-15 AS=76.8e-15 PD=1.26e-6 PS=1.26e-6 NRD=1.16667 NRS=1.16667 M=1
mi14__i16__pm9 n406__vdd i14__i16__net5 n10__i14__i16__net4 n293__vdd g45p1svt L=45e-9 W=480e-9 AD=67.2e-15 AS=67.2e-15 PD=1.26e-6 PS=1.26e-6 NRD=1.16667 NRS=1.16667 M=1
mi14__i16__pm11 n10__i14__y_out_b_0 n4__i14__i16__net4 n404__vdd n293__vdd g45p1svt L=45e-9 W=480e-9 AD=67.2e-15 AS=67.2e-15 PD=1.24e-6 PS=1.24e-6 NRD=1.16667 NRS=1.16667 M=1
mi14__i16__pm13 x_out_2 i14__y_out_b_0 n402__vdd n293__vdd g45p1svt L=45e-9 W=480e-9 AD=67.2e-15 AS=67.2e-15 PD=1.24e-6 PS=1.24e-6 NRD=1.16667 NRS=1.16667 M=1
mi14__i12__pm0 n13__i14__i12__net1 n36__i14__net10 n1__y0 n32__vdd g45p1svt L=45e-9 W=120e-9 AD=16.8e-15 AS=16.8e-15 PD=520e-9 PS=520e-9 NRD=1.16667 NRS=1.16667 M=1
mi14__i12__pm2 n105__vdd n3__i14__i12__net2 n9__i14__i12__net1 n32__vdd g45p1svt L=180e-9 W=120e-9 AD=16.8e-15 AS=16.8e-15 PD=520e-9 PS=520e-9 NRD=1.16667 NRS=1.16667 M=1
mi14__i12__pm1_1__rcx n11__i14__i12__net2 n7__i14__i12__net1 n103__vdd n32__vdd g45p1svt L=45e-9 W=480e-9 AD=76.8e-15 AS=76.8e-15 PD=1.26e-6 PS=1.26e-6 NRD=1.16667 NRS=1.16667 M=1
mi14__i12__pm1 n101__vdd i14__i12__net1 n11__i14__i12__net2 n32__vdd g45p1svt L=45e-9 W=480e-9 AD=67.2e-15 AS=67.2e-15 PD=1.26e-6 PS=1.26e-6 NRD=1.16667 NRS=1.16667 M=1
mi14__i12__pm8 n13__i14__i12__net5 n56__i14__net9 n6__i14__i12__net2 n32__vdd g45p1svt L=45e-9 W=120e-9 AD=16.8e-15 AS=16.8e-15 PD=520e-9 PS=520e-9 NRD=1.16667 NRS=1.16667 M=1
mi14__i12__pm10 n99__vdd n3__i14__i12__net4 n9__i14__i12__net5 n32__vdd g45p1svt L=180e-9 W=120e-9 AD=16.8e-15 AS=16.8e-15 PD=520e-9 PS=520e-9 NRD=1.16667 NRS=1.16667 M=1
mi14__i12__pm15 n15__i14__i12__net5 n27__i14__net4 n97__vdd n32__vdd g45p1svt L=45e-9 W=120e-9 AD=16.8e-15 AS=16.8e-15 PD=520e-9 PS=520e-9 NRD=1.16667 NRS=1.16667 M=1
mi14__i12__pm9_1__rcx n11__i14__i12__net4 n7__i14__i12__net5 n95__vdd n32__vdd g45p1svt L=45e-9 W=480e-9 AD=76.8e-15 AS=76.8e-15 PD=1.26e-6 PS=1.26e-6 NRD=1.16667 NRS=1.16667 M=1
mi14__i12__pm9 n93__vdd i14__i12__net5 n11__i14__i12__net4 n32__vdd g45p1svt L=45e-9 W=480e-9 AD=67.2e-15 AS=67.2e-15 PD=1.26e-6 PS=1.26e-6 NRD=1.16667 NRS=1.16667 M=1
mi14__i12__pm11 n10__i14__x_out_b_0 n4__i14__i12__net4 n91__vdd n32__vdd g45p1svt L=45e-9 W=480e-9 AD=67.2e-15 AS=67.2e-15 PD=1.24e-6 PS=1.24e-6 NRD=1.16667 NRS=1.16667 M=1
mi14__i12__pm13 n9__y_out_0 i14__x_out_b_0 n89__vdd n32__vdd g45p1svt L=45e-9 W=480e-9 AD=67.2e-15 AS=67.2e-15 PD=1.24e-6 PS=1.24e-6 NRD=1.16667 NRS=1.16667 M=1
mi14__i9__pm0 n13__i14__i9__net1 n8__i14__net10 n1__x0 n32__vdd g45p1svt L=45e-9 W=120e-9 AD=16.8e-15 AS=16.8e-15 PD=520e-9 PS=520e-9 NRD=1.16667 NRS=1.16667 M=1
mi14__i9__pm2 n126__vdd n3__i14__i9__net2 n9__i14__i9__net1 n32__vdd g45p1svt L=180e-9 W=120e-9 AD=16.8e-15 AS=16.8e-15 PD=520e-9 PS=520e-9 NRD=1.16667 NRS=1.16667 M=1
mi14__i9__pm1_1__rcx n11__i14__i9__net2 n7__i14__i9__net1 n122__vdd n32__vdd g45p1svt L=45e-9 W=480e-9 AD=76.8e-15 AS=76.8e-15 PD=1.26e-6 PS=1.26e-6 NRD=1.16667 NRS=1.16667 M=1
mi14__i9__pm1 n119__vdd i14__i9__net1 n11__i14__i9__net2 n32__vdd g45p1svt L=45e-9 W=480e-9 AD=67.2e-15 AS=67.2e-15 PD=1.26e-6 PS=1.26e-6 NRD=1.16667 NRS=1.16667 M=1
mi14__i9__pm8 n13__i14__i9__net5 n16__i14__net9 n6__i14__i9__net2 n32__vdd g45p1svt L=45e-9 W=120e-9 AD=16.8e-15 AS=16.8e-15 PD=520e-9 PS=520e-9 NRD=1.16667 NRS=1.16667 M=1
mi14__i9__pm10 n117__vdd n3__i14__i9__net4 n9__i14__i9__net5 n32__vdd g45p1svt L=180e-9 W=120e-9 AD=16.8e-15 AS=16.8e-15 PD=520e-9 PS=520e-9 NRD=1.16667 NRS=1.16667 M=1
mi14__i9__pm15 n15__i14__i9__net5 n7__i14__net4 n115__vdd n32__vdd g45p1svt L=45e-9 W=120e-9 AD=16.8e-15 AS=16.8e-15 PD=520e-9 PS=520e-9 NRD=1.16667 NRS=1.16667 M=1
mi14__i9__pm9_1__rcx n10__i14__i9__net4 n7__i14__i9__net5 n113__vdd n32__vdd g45p1svt L=45e-9 W=480e-9 AD=76.8e-15 AS=76.8e-15 PD=1.26e-6 PS=1.26e-6 NRD=1.16667 NRS=1.16667 M=1
mi14__i9__pm9 n111__vdd i14__i9__net5 n10__i14__i9__net4 n32__vdd g45p1svt L=45e-9 W=480e-9 AD=67.2e-15 AS=67.2e-15 PD=1.26e-6 PS=1.26e-6 NRD=1.16667 NRS=1.16667 M=1
mi14__i9__pm11 n10__i14__x_out_b_3 n4__i14__i9__net4 n109__vdd n32__vdd g45p1svt L=45e-9 W=480e-9 AD=67.2e-15 AS=67.2e-15 PD=1.24e-6 PS=1.24e-6 NRD=1.16667 NRS=1.16667 M=1
mi14__i9__pm13 x_out_0 i14__x_out_b_3 n107__vdd n32__vdd g45p1svt L=45e-9 W=480e-9 AD=67.2e-15 AS=67.2e-15 PD=1.24e-6 PS=1.24e-6 NRD=1.16667 NRS=1.16667 M=1
mi14__pm9 n2__ck4 n4__i14__net11 n253__vdd n134__vdd g45p1svt L=45e-9 W=480e-9 AD=67.2e-15 AS=67.2e-15 PD=1.24e-6 PS=1.24e-6 NRD=1.16667 NRS=1.16667 M=1
mi14__pm10 i14__clk_div4_out_b n4__i14__net7 n255__vdd n134__vdd g45p1svt L=45e-9 W=480e-9 AD=67.2e-15 AS=67.2e-15 PD=1.24e-6 PS=1.24e-6 NRD=1.16667 NRS=1.16667 M=1
mi13__i20__i4__pm2 n5__i13__i20__i4__net2 n8__i13__net18 n68__vdd n32__vdd g45p1svt L=45e-9 W=240e-9 AD=33.6e-15 AS=33.6e-15 PD=760e-9 PS=760e-9 NRD=1.16667 NRS=1.16667 M=1
mi13__i20__i4__pm0 n6__r1 n9__i13__net18 n18__i13__net7 n32__vdd g45p1svt L=45e-9 W=120e-9 AD=16.8e-15 AS=16.8e-15 PD=520e-9 PS=520e-9 NRD=1.16667 NRS=1.16667 M=1
mi13__i20__i4__pm1 n10__r1 n8__i13__net7 n26__i13__net18 n32__vdd g45p1svt L=45e-9 W=240e-9 AD=33.6e-15 AS=33.6e-15 PD=760e-9 PS=760e-9 NRD=1.16667 NRS=1.16667 M=1
mi13__i20__pm0 n10__i13__i20__net1 n4__i13__net18 n71__vdd n32__vdd g45p1svt L=45e-9 W=240e-9 AD=33.6e-15 AS=33.6e-15 PD=780e-9 PS=780e-9 NRD=1.16667 NRS=1.16667 M=1
mi13__i20__pm1 n71__vdd n4__i13__net7 n6__i13__i20__net1 n32__vdd g45p1svt L=45e-9 W=240e-9 AD=38.4e-15 AS=38.4e-15 PD=780e-9 PS=780e-9 NRD=1.16667 NRS=1.16667 M=1
mi13__i20__pm2 n9__i13__net23 n4__i13__i20__net1 n70__vdd n32__vdd g45p1svt L=45e-9 W=240e-9 AD=33.6e-15 AS=33.6e-15 PD=760e-9 PS=760e-9 NRD=1.16667 NRS=1.16667 M=1
mi13__i19__i4__pm2 n5__i13__i19__i4__net2 n8__i13__net1 n74__vdd n32__vdd g45p1svt L=45e-9 W=240e-9 AD=33.6e-15 AS=33.6e-15 PD=760e-9 PS=760e-9 NRD=1.16667 NRS=1.16667 M=1
mi13__i19__i4__pm0 n12__i13__net18 n9__i13__net1 n18__i13__net11 n32__vdd g45p1svt L=45e-9 W=120e-9 AD=16.8e-15 AS=16.8e-15 PD=520e-9 PS=520e-9 NRD=1.16667 NRS=1.16667 M=1
mi13__i19__i4__pm1 n16__i13__net18 n8__i13__net11 n22__i13__net1 n32__vdd g45p1svt L=45e-9 W=240e-9 AD=33.6e-15 AS=33.6e-15 PD=760e-9 PS=760e-9 NRD=1.16667 NRS=1.16667 M=1
mi13__i19__pm0 n10__i13__i19__net1 n4__i13__net1 n78__vdd n32__vdd g45p1svt L=45e-9 W=240e-9 AD=33.6e-15 AS=33.6e-15 PD=780e-9 PS=780e-9 NRD=1.16667 NRS=1.16667 M=1
mi13__i19__pm1 n78__vdd n4__i13__net11 n6__i13__i19__net1 n32__vdd g45p1svt L=45e-9 W=240e-9 AD=38.4e-15 AS=38.4e-15 PD=780e-9 PS=780e-9 NRD=1.16667 NRS=1.16667 M=1
mi13__i19__pm2 n8__i13__net17 n4__i13__i19__net1 n76__vdd n32__vdd g45p1svt L=45e-9 W=240e-9 AD=33.6e-15 AS=33.6e-15 PD=760e-9 PS=760e-9 NRD=1.16667 NRS=1.16667 M=1
mi13__i17__i4__pm2 n5__i13__i17__i4__net2 n8__i13__a2 n80__vdd n32__vdd g45p1svt L=45e-9 W=240e-9 AD=33.6e-15 AS=33.6e-15 PD=760e-9 PS=760e-9 NRD=1.16667 NRS=1.16667 M=1
mi13__i17__i4__pm0 n10__i13__net12 n13__i13__a2 n22__i13__a3 n32__vdd g45p1svt L=45e-9 W=120e-9 AD=16.8e-15 AS=16.8e-15 PD=520e-9 PS=520e-9 NRD=1.16667 NRS=1.16667 M=1
mi13__i17__i4__pm1 n14__i13__net12 n8__i13__a3 n28__i13__a2 n32__vdd g45p1svt L=45e-9 W=240e-9 AD=33.6e-15 AS=33.6e-15 PD=760e-9 PS=760e-9 NRD=1.16667 NRS=1.16667 M=1
mi13__i17__pm0 n10__i13__i17__net1 n4__i13__a2 n84__vdd n32__vdd g45p1svt L=45e-9 W=240e-9 AD=33.6e-15 AS=33.6e-15 PD=780e-9 PS=780e-9 NRD=1.16667 NRS=1.16667 M=1
mi13__i17__pm1 n84__vdd n4__i13__a3 n6__i13__i17__net1 n32__vdd g45p1svt L=45e-9 W=240e-9 AD=38.4e-15 AS=38.4e-15 PD=780e-9 PS=780e-9 NRD=1.16667 NRS=1.16667 M=1
mi13__i17__pm2 n12__i13__net11 n4__i13__i17__net1 n82__vdd n32__vdd g45p1svt L=45e-9 W=240e-9 AD=33.6e-15 AS=33.6e-15 PD=760e-9 PS=760e-9 NRD=1.16667 NRS=1.16667 M=1
mi13__i18__i4__pm2 n3__i13__i18__i4__net2 n5__i13__net2 n73__vdd n32__vdd g45p1svt L=45e-9 W=240e-9 AD=33.6e-15 AS=33.6e-15 PD=760e-9 PS=760e-9 NRD=1.16667 NRS=1.16667 M=1
mi13__i18__i4__pm0 n2__r0 n9__i13__net2 n22__i13__net12 n32__vdd g45p1svt L=45e-9 W=120e-9 AD=16.8e-15 AS=16.8e-15 PD=520e-9 PS=520e-9 NRD=1.16667 NRS=1.16667 M=1
mi13__i18__i4__pm1 n5__r0 n5__i13__net12 n26__i13__net2 n32__vdd g45p1svt L=45e-9 W=240e-9 AD=33.6e-15 AS=33.6e-15 PD=760e-9 PS=760e-9 NRD=1.16667 NRS=1.16667 M=1
mi13__i18__pm0 n10__i13__i18__net1 i13__net2 n77__vdd n32__vdd g45p1svt L=45e-9 W=240e-9 AD=33.6e-15 AS=33.6e-15 PD=780e-9 PS=780e-9 NRD=1.16667 NRS=1.16667 M=1
mi13__i18__pm1 n77__vdd i13__net12 n5__i13__i18__net1 n32__vdd g45p1svt L=45e-9 W=240e-9 AD=38.4e-15 AS=38.4e-15 PD=780e-9 PS=780e-9 NRD=1.16667 NRS=1.16667 M=1
mi13__i18__pm2 n12__i13__net7 i13__i18__net1 n75__vdd n32__vdd g45p1svt L=45e-9 W=240e-9 AD=33.6e-15 AS=33.6e-15 PD=760e-9 PS=760e-9 NRD=1.16667 NRS=1.16667 M=1
mi13__i16__i4__pm2 n3__i13__i16__i4__net2 n5__i13__a0 n79__vdd n32__vdd g45p1svt L=45e-9 W=240e-9 AD=33.6e-15 AS=33.6e-15 PD=760e-9 PS=760e-9 NRD=1.16667 NRS=1.16667 M=1
mi13__i16__i4__pm0 n12__i13__net2 n13__i13__a0 n22__i13__a1 n32__vdd g45p1svt L=45e-9 W=120e-9 AD=16.8e-15 AS=16.8e-15 PD=520e-9 PS=520e-9 NRD=1.16667 NRS=1.16667 M=1
mi13__i16__i4__pm1 n15__i13__net2 n5__i13__a1 n28__i13__a0 n32__vdd g45p1svt L=45e-9 W=240e-9 AD=33.6e-15 AS=33.6e-15 PD=760e-9 PS=760e-9 NRD=1.16667 NRS=1.16667 M=1
mi13__i16__pm0 n10__i13__i16__net1 i13__a0 n83__vdd n32__vdd g45p1svt L=45e-9 W=240e-9 AD=33.6e-15 AS=33.6e-15 PD=780e-9 PS=780e-9 NRD=1.16667 NRS=1.16667 M=1
mi13__i16__pm1 n83__vdd i13__a1 n5__i13__i16__net1 n32__vdd g45p1svt L=45e-9 W=240e-9 AD=38.4e-15 AS=38.4e-15 PD=780e-9 PS=780e-9 NRD=1.16667 NRS=1.16667 M=1
mi13__i16__pm2 n14__i13__net1 i13__i16__net1 n81__vdd n32__vdd g45p1svt L=45e-9 W=240e-9 AD=33.6e-15 AS=33.6e-15 PD=760e-9 PS=760e-9 NRD=1.16667 NRS=1.16667 M=1
mi13__i15__pm2 n5__i13__i15__net2 n9__x_out_3 n86__vdd n32__vdd g45p1svt L=45e-9 W=240e-9 AD=33.6e-15 AS=33.6e-15 PD=760e-9 PS=760e-9 NRD=1.16667 NRS=1.16667 M=1
mi13__i15__pm0 n10__i13__a3 n10__x_out_3 n15__y_out_3 n32__vdd g45p1svt L=45e-9 W=120e-9 AD=16.8e-15 AS=16.8e-15 PD=520e-9 PS=520e-9 NRD=1.16667 NRS=1.16667 M=1
mi13__i15__pm1 n14__i13__a3 n4__y_out_3 n21__x_out_3 n32__vdd g45p1svt L=45e-9 W=240e-9 AD=33.6e-15 AS=33.6e-15 PD=760e-9 PS=760e-9 NRD=1.16667 NRS=1.16667 M=1
mi13__i14__pm2 n5__i13__i14__net2 n9__x_out_2 n88__vdd n32__vdd g45p1svt L=45e-9 W=240e-9 AD=33.6e-15 AS=33.6e-15 PD=760e-9 PS=760e-9 NRD=1.16667 NRS=1.16667 M=1
mi13__i14__pm0 n10__i13__a2 n10__x_out_2 n14__y_out_2 n32__vdd g45p1svt L=45e-9 W=120e-9 AD=16.8e-15 AS=16.8e-15 PD=520e-9 PS=520e-9 NRD=1.16667 NRS=1.16667 M=1
mi13__i14__pm1 n16__i13__a2 n4__y_out_2 n22__x_out_2 n32__vdd g45p1svt L=45e-9 W=240e-9 AD=33.6e-15 AS=33.6e-15 PD=760e-9 PS=760e-9 NRD=1.16667 NRS=1.16667 M=1
mi13__i13__pm2 n3__i13__i13__net2 n6__x_out_1 n85__vdd n32__vdd g45p1svt L=45e-9 W=240e-9 AD=33.6e-15 AS=33.6e-15 PD=760e-9 PS=760e-9 NRD=1.16667 NRS=1.16667 M=1
mi13__i13__pm0 n10__i13__a1 n10__x_out_1 n14__y_out_1 n32__vdd g45p1svt L=45e-9 W=120e-9 AD=16.8e-15 AS=16.8e-15 PD=520e-9 PS=520e-9 NRD=1.16667 NRS=1.16667 M=1
mi13__i13__pm1 n13__i13__a1 y_out_1 n22__x_out_1 n32__vdd g45p1svt L=45e-9 W=240e-9 AD=33.6e-15 AS=33.6e-15 PD=760e-9 PS=760e-9 NRD=1.16667 NRS=1.16667 M=1
mi13__i12__pm2 n3__i13__i12__net2 y_out_0 n87__vdd n32__vdd g45p1svt L=45e-9 W=240e-9 AD=33.6e-15 AS=33.6e-15 PD=760e-9 PS=760e-9 NRD=1.16667 NRS=1.16667 M=1
mi13__i12__pm0 n10__i13__a0 n5__y_out_0 n16__x_out_0 n32__vdd g45p1svt L=45e-9 W=120e-9 AD=16.8e-15 AS=16.8e-15 PD=520e-9 PS=520e-9 NRD=1.16667 NRS=1.16667 M=1
mi13__i12__pm1 n15__i13__a0 n6__x_out_0 n18__y_out_0 n32__vdd g45p1svt L=45e-9 W=240e-9 AD=33.6e-15 AS=33.6e-15 PD=760e-9 PS=760e-9 NRD=1.16667 NRS=1.16667 M=1
mi13__pm0 n7__i13__net3 i13__net23 i13__net6 n32__vdd g45p1svt L=45e-9 W=480e-9 AD=67.2e-15 AS=67.2e-15 PD=1.26e-6 PS=1.26e-6 NRD=1.16667 NRS=1.16667 M=1
mi13__pm1 i13__net6 i13__net17 n72__vdd n32__vdd g45p1svt L=45e-9 W=480e-9 AD=76.8e-15 AS=76.8e-15 PD=1.26e-6 PS=1.26e-6 NRD=1.16667 NRS=1.16667 M=1
mi13__pm2 r2 i13__net3 n69__vdd n32__vdd g45p1svt L=45e-9 W=240e-9 AD=33.6e-15 AS=33.6e-15 PD=760e-9 PS=760e-9 NRD=1.16667 NRS=1.16667 M=1
mi9__i1__pm1_1__rcx n25__shift n6__i9__net1 n226__vdd n134__vdd g45p1svt L=45e-9 W=360e-9 AD=57.6e-15 AS=57.6e-15 PD=1.02e-6 PS=1.02e-6 NRD=1.16667 NRS=1.16667 M=1
mi9__i1__pm1 n225__vdd i9__net1 n25__shift n134__vdd g45p1svt L=45e-9 W=360e-9 AD=57.6e-15 AS=57.6e-15 PD=1.04e-6 PS=1.04e-6 NRD=1.16667 NRS=1.16667 M=1
mi9__i1__pm0_1__rcx n29__shift n15__ck4 n225__vdd n134__vdd g45p1svt L=45e-9 W=360e-9 AD=57.6e-15 AS=57.6e-15 PD=1.04e-6 PS=1.04e-6 NRD=1.16667 NRS=1.16667 M=1
mi9__i1__pm0 n224__vdd n10__ck4 n29__shift n134__vdd g45p1svt L=45e-9 W=360e-9 AD=50.4e-15 AS=50.4e-15 PD=1.02e-6 PS=1.02e-6 NRD=1.16667 NRS=1.16667 M=1
mi9__i4__pm0 n13__i9__i4__net1 n2__ck_buff n6__ck4 n134__vdd g45p1svt L=45e-9 W=120e-9 AD=16.8e-15 AS=16.8e-15 PD=520e-9 PS=520e-9 NRD=1.16667 NRS=1.16667 M=1
mi9__i4__pm2 n241__vdd n3__i9__i4__net2 n9__i9__i4__net1 n134__vdd g45p1svt L=180e-9 W=120e-9 AD=16.8e-15 AS=16.8e-15 PD=520e-9 PS=520e-9 NRD=1.16667 NRS=1.16667 M=1
mi9__i4__pm1_1__rcx n11__i9__i4__net2 n7__i9__i4__net1 n238__vdd n134__vdd g45p1svt L=45e-9 W=480e-9 AD=76.8e-15 AS=76.8e-15 PD=1.26e-6 PS=1.26e-6 NRD=1.16667 NRS=1.16667 M=1
mi9__i4__pm1 n236__vdd i9__i4__net1 n11__i9__i4__net2 n134__vdd g45p1svt L=45e-9 W=480e-9 AD=67.2e-15 AS=67.2e-15 PD=1.26e-6 PS=1.26e-6 NRD=1.16667 NRS=1.16667 M=1
mi9__i4__pm8 n13__i9__i4__net5 n4__ck_b n6__i9__i4__net2 n134__vdd g45p1svt L=45e-9 W=120e-9 AD=16.8e-15 AS=16.8e-15 PD=520e-9 PS=520e-9 NRD=1.16667 NRS=1.16667 M=1
mi9__i4__pm10 n235__vdd n3__i9__i4__net4 n9__i9__i4__net5 n134__vdd g45p1svt L=180e-9 W=120e-9 AD=16.8e-15 AS=16.8e-15 PD=520e-9 PS=520e-9 NRD=1.16667 NRS=1.16667 M=1
mi9__i4__pm15 n15__i9__i4__net5 reset_b n234__vdd n134__vdd g45p1svt L=45e-9 W=120e-9 AD=16.8e-15 AS=16.8e-15 PD=520e-9 PS=520e-9 NRD=1.16667 NRS=1.16667 M=1
mi9__i4__pm9_1__rcx n10__i9__i4__net4 n7__i9__i4__net5 n233__vdd n134__vdd g45p1svt L=45e-9 W=480e-9 AD=76.8e-15 AS=76.8e-15 PD=1.26e-6 PS=1.26e-6 NRD=1.16667 NRS=1.16667 M=1
mi9__i4__pm9 n231__vdd i9__i4__net5 n10__i9__i4__net4 n134__vdd g45p1svt L=45e-9 W=480e-9 AD=67.2e-15 AS=67.2e-15 PD=1.26e-6 PS=1.26e-6 NRD=1.16667 NRS=1.16667 M=1
mi9__i4__pm11 n8__i9__net2 n4__i9__i4__net4 n229__vdd n134__vdd g45p1svt L=45e-9 W=480e-9 AD=67.2e-15 AS=67.2e-15 PD=1.24e-6 PS=1.24e-6 NRD=1.16667 NRS=1.16667 M=1
mi9__i4__pm13 n7__i9__net1 i9__net2 n227__vdd n134__vdd g45p1svt L=45e-9 W=480e-9 AD=67.2e-15 AS=67.2e-15 PD=1.24e-6 PS=1.24e-6 NRD=1.16667 NRS=1.16667 M=1
mi12__pm0 n14__i12__bcore_bar n13__serial_out n130__vdd n132__vdd g45p1svt L=45e-9 W=240e-9 AD=33.6e-15 AS=33.6e-15 PD=760e-9 PS=760e-9 NRD=1.16667 NRS=1.16667 M=1
mi40__m0 n6__serial_out_b_high_buff n4__serial_out_b_high n1010__vss n640__vss g45n2svt L=150e-9 W=320e-9 AD=48e-15 AS=48e-15 PD=940e-9 PS=940e-9 NRD=468.75e-3 NRS=468.75e-3 M=1
mi18__m15_99__rcx n31__r_out n16__i18__net5 n1284__vss n640__vss g45n2svt L=150e-9 W=6e-6 AD=1.2e-12 AS=1.2e-12 PD=12.4e-6 PS=12.4e-6 NRD=468.75e-3 NRS=468.75e-3 M=1
mi18__m15_98__rcx n1288__vss n13__i18__net5 n31__r_out n640__vss g45n2svt L=150e-9 W=6e-6 AD=1.2e-12 AS=1.2e-12 PD=12.4e-6 PS=12.4e-6 NRD=468.75e-3 NRS=468.75e-3 M=1
mi18__m15_97__rcx n14__r_out n10__i18__net5 n1288__vss n640__vss g45n2svt L=150e-9 W=6e-6 AD=1.2e-12 AS=1.2e-12 PD=12.4e-6 PS=12.4e-6 NRD=468.75e-3 NRS=468.75e-3 M=1
mi18__m15_96__rcx n1292__vss n7__i18__net5 n14__r_out n640__vss g45n2svt L=150e-9 W=6e-6 AD=1.2e-12 AS=1.2e-12 PD=12.4e-6 PS=12.4e-6 NRD=468.75e-3 NRS=468.75e-3 M=1
mi18__m15_95__rcx n7__r_out n4__i18__net5 n1292__vss n640__vss g45n2svt L=150e-9 W=6e-6 AD=1.2e-12 AS=1.2e-12 PD=12.4e-6 PS=12.4e-6 NRD=468.75e-3 NRS=468.75e-3 M=1
mi18__m15_94__rcx n1295__vss i18__net5 n7__r_out n640__vss g45n2svt L=150e-9 W=6e-6 AD=900e-15 AS=900e-15 PD=12.35e-6 PS=12.35e-6 NRD=468.75e-3 NRS=468.75e-3 M=1
mi18__m15_93__rcx n72__r_out n34__i18__net5 n1272__vss n640__vss g45n2svt L=150e-9 W=6e-6 AD=1.2e-12 AS=1.2e-12 PD=12.4e-6 PS=12.4e-6 NRD=468.75e-3 NRS=468.75e-3 M=1
mi18__m15_92__rcx n1276__vss n31__i18__net5 n72__r_out n640__vss g45n2svt L=150e-9 W=6e-6 AD=1.2e-12 AS=1.2e-12 PD=12.4e-6 PS=12.4e-6 NRD=468.75e-3 NRS=468.75e-3 M=1
mi18__m15_91__rcx n57__r_out n28__i18__net5 n1276__vss n640__vss g45n2svt L=150e-9 W=6e-6 AD=1.2e-12 AS=1.2e-12 PD=12.4e-6 PS=12.4e-6 NRD=468.75e-3 NRS=468.75e-3 M=1
mi18__m15_90__rcx n1280__vss n25__i18__net5 n57__r_out n640__vss g45n2svt L=150e-9 W=6e-6 AD=1.2e-12 AS=1.2e-12 PD=12.4e-6 PS=12.4e-6 NRD=468.75e-3 NRS=468.75e-3 M=1
mi18__m15_89__rcx n46__r_out n22__i18__net5 n1280__vss n640__vss g45n2svt L=150e-9 W=6e-6 AD=1.2e-12 AS=1.2e-12 PD=12.4e-6 PS=12.4e-6 NRD=468.75e-3 NRS=468.75e-3 M=1
mi18__m15_88__rcx n1284__vss n19__i18__net5 n46__r_out n640__vss g45n2svt L=150e-9 W=6e-6 AD=1.2e-12 AS=1.2e-12 PD=12.4e-6 PS=12.4e-6 NRD=468.75e-3 NRS=468.75e-3 M=1
mi18__m15_87__rcx n1272__vss n37__i18__net5 n79__r_out n640__vss g45n2svt L=150e-9 W=6e-6 AD=1.2e-12 AS=1.2e-12 PD=12.4e-6 PS=12.4e-6 NRD=468.75e-3 NRS=468.75e-3 M=1
mi18__m15_86__rcx n1259__vss n63__i18__net5 n124__r_out n640__vss g45n2svt L=150e-9 W=6e-6 AD=1.2e-12 AS=1.2e-12 PD=12.4e-6 PS=12.4e-6 NRD=468.75e-3 NRS=468.75e-3 M=1
mi18__m15_85__rcx n111__r_out n60__i18__net5 n1259__vss n640__vss g45n2svt L=150e-9 W=6e-6 AD=1.2e-12 AS=1.2e-12 PD=12.4e-6 PS=12.4e-6 NRD=468.75e-3 NRS=468.75e-3 M=1
mi18__m15_84__rcx n1263__vss n53__i18__net5 n111__r_out n640__vss g45n2svt L=150e-9 W=6e-6 AD=1.2e-12 AS=1.2e-12 PD=12.4e-6 PS=12.4e-6 NRD=468.75e-3 NRS=468.75e-3 M=1
mi18__m15_83__rcx n98__r_out n50__i18__net5 n1263__vss n640__vss g45n2svt L=150e-9 W=6e-6 AD=1.2e-12 AS=1.2e-12 PD=12.4e-6 PS=12.4e-6 NRD=468.75e-3 NRS=468.75e-3 M=1
mi18__m15_82__rcx n1268__vss n43__i18__net5 n98__r_out n640__vss g45n2svt L=150e-9 W=6e-6 AD=1.2e-12 AS=1.2e-12 PD=12.4e-6 PS=12.4e-6 NRD=468.75e-3 NRS=468.75e-3 M=1
mi18__m15_81__rcx n79__r_out n40__i18__net5 n1268__vss n640__vss g45n2svt L=150e-9 W=6e-6 AD=1.2e-12 AS=1.2e-12 PD=12.4e-6 PS=12.4e-6 NRD=468.75e-3 NRS=468.75e-3 M=1
mi18__m15_80__rcx n1247__vss n95__i18__net5 n161__r_out n640__vss g45n2svt L=150e-9 W=6e-6 AD=1.2e-12 AS=1.2e-12 PD=12.4e-6 PS=12.4e-6 NRD=468.75e-3 NRS=468.75e-3 M=1
mi18__m15_79__rcx n144__r_out n90__i18__net5 n1247__vss n640__vss g45n2svt L=150e-9 W=6e-6 AD=1.2e-12 AS=1.2e-12 PD=12.4e-6 PS=12.4e-6 NRD=468.75e-3 NRS=468.75e-3 M=1
mi18__m15_78__rcx n1251__vss n85__i18__net5 n144__r_out n640__vss g45n2svt L=150e-9 W=6e-6 AD=1.2e-12 AS=1.2e-12 PD=12.4e-6 PS=12.4e-6 NRD=468.75e-3 NRS=468.75e-3 M=1
mi18__m15_77__rcx n131__r_out n78__i18__net5 n1251__vss n640__vss g45n2svt L=150e-9 W=6e-6 AD=1.2e-12 AS=1.2e-12 PD=12.4e-6 PS=12.4e-6 NRD=468.75e-3 NRS=468.75e-3 M=1
mi18__m15_76__rcx n1255__vss n73__i18__net5 n131__r_out n640__vss g45n2svt L=150e-9 W=6e-6 AD=1.2e-12 AS=1.2e-12 PD=12.4e-6 PS=12.4e-6 NRD=468.75e-3 NRS=468.75e-3 M=1
mi18__m15_75__rcx n124__r_out n68__i18__net5 n1255__vss n640__vss g45n2svt L=150e-9 W=6e-6 AD=1.2e-12 AS=1.2e-12 PD=12.4e-6 PS=12.4e-6 NRD=468.75e-3 NRS=468.75e-3 M=1
mi18__m15_74__rcx n1234__vss n123__i18__net5 n202__r_out n640__vss g45n2svt L=150e-9 W=6e-6 AD=1.2e-12 AS=1.2e-12 PD=12.4e-6 PS=12.4e-6 NRD=468.75e-3 NRS=468.75e-3 M=1
mi18__m15_73__rcx n187__r_out n120__i18__net5 n1234__vss n640__vss g45n2svt L=150e-9 W=6e-6 AD=1.2e-12 AS=1.2e-12 PD=12.4e-6 PS=12.4e-6 NRD=468.75e-3 NRS=468.75e-3 M=1
mi18__m15_72__rcx n1239__vss n115__i18__net5 n187__r_out n640__vss g45n2svt L=150e-9 W=6e-6 AD=1.2e-12 AS=1.2e-12 PD=12.4e-6 PS=12.4e-6 NRD=468.75e-3 NRS=468.75e-3 M=1
mi18__m15_71__rcx n176__r_out n110__i18__net5 n1239__vss n640__vss g45n2svt L=150e-9 W=6e-6 AD=1.2e-12 AS=1.2e-12 PD=12.4e-6 PS=12.4e-6 NRD=468.75e-3 NRS=468.75e-3 M=1
mi18__m15_70__rcx n1243__vss n103__i18__net5 n176__r_out n640__vss g45n2svt L=150e-9 W=6e-6 AD=1.2e-12 AS=1.2e-12 PD=12.4e-6 PS=12.4e-6 NRD=468.75e-3 NRS=468.75e-3 M=1
mi18__m15_69__rcx n161__r_out n100__i18__net5 n1243__vss n640__vss g45n2svt L=150e-9 W=6e-6 AD=1.2e-12 AS=1.2e-12 PD=12.4e-6 PS=12.4e-6 NRD=468.75e-3 NRS=468.75e-3 M=1
mi18__m15_68__rcx n1221__vss n153__i18__net5 n241__r_out n640__vss g45n2svt L=150e-9 W=6e-6 AD=1.2e-12 AS=1.2e-12 PD=12.4e-6 PS=12.4e-6 NRD=468.75e-3 NRS=468.75e-3 M=1
mi18__m15_67__rcx n228__r_out n148__i18__net5 n1221__vss n640__vss g45n2svt L=150e-9 W=6e-6 AD=1.2e-12 AS=1.2e-12 PD=12.4e-6 PS=12.4e-6 NRD=468.75e-3 NRS=468.75e-3 M=1
mi18__m15_66__rcx n1226__vss n143__i18__net5 n228__r_out n640__vss g45n2svt L=150e-9 W=6e-6 AD=1.2e-12 AS=1.2e-12 PD=12.4e-6 PS=12.4e-6 NRD=468.75e-3 NRS=468.75e-3 M=1
mi18__m15_65__rcx n209__r_out n138__i18__net5 n1226__vss n640__vss g45n2svt L=150e-9 W=6e-6 AD=1.2e-12 AS=1.2e-12 PD=12.4e-6 PS=12.4e-6 NRD=468.75e-3 NRS=468.75e-3 M=1
mi18__m15_64__rcx n1230__vss n135__i18__net5 n209__r_out n640__vss g45n2svt L=150e-9 W=6e-6 AD=1.2e-12 AS=1.2e-12 PD=12.4e-6 PS=12.4e-6 NRD=468.75e-3 NRS=468.75e-3 M=1
mi18__m15_63__rcx n202__r_out n129__i18__net5 n1230__vss n640__vss g45n2svt L=150e-9 W=6e-6 AD=1.2e-12 AS=1.2e-12 PD=12.4e-6 PS=12.4e-6 NRD=468.75e-3 NRS=468.75e-3 M=1
mi18__m15_62__rcx n241__r_out n160__i18__net5 n1217__vss n640__vss g45n2svt L=150e-9 W=6e-6 AD=1.2e-12 AS=1.2e-12 PD=12.4e-6 PS=12.4e-6 NRD=468.75e-3 NRS=468.75e-3 M=1
mi18__m15_61__rcx n274__r_out n188__i18__net5 n1204__vss n640__vss g45n2svt L=150e-9 W=6e-6 AD=1.2e-12 AS=1.2e-12 PD=12.4e-6 PS=12.4e-6 NRD=468.75e-3 NRS=468.75e-3 M=1
mi18__m15_60__rcx n1209__vss n185__i18__net5 n274__r_out n640__vss g45n2svt L=150e-9 W=6e-6 AD=1.2e-12 AS=1.2e-12 PD=12.4e-6 PS=12.4e-6 NRD=468.75e-3 NRS=468.75e-3 M=1
mi18__m15_59__rcx n267__r_out n179__i18__net5 n1209__vss n640__vss g45n2svt L=150e-9 W=6e-6 AD=1.2e-12 AS=1.2e-12 PD=12.4e-6 PS=12.4e-6 NRD=468.75e-3 NRS=468.75e-3 M=1
mi18__m15_58__rcx n1213__vss n173__i18__net5 n267__r_out n640__vss g45n2svt L=150e-9 W=6e-6 AD=1.2e-12 AS=1.2e-12 PD=12.4e-6 PS=12.4e-6 NRD=468.75e-3 NRS=468.75e-3 M=1
mi18__m15_57__rcx n254__r_out n170__i18__net5 n1213__vss n640__vss g45n2svt L=150e-9 W=6e-6 AD=1.2e-12 AS=1.2e-12 PD=12.4e-6 PS=12.4e-6 NRD=468.75e-3 NRS=468.75e-3 M=1
mi18__m15_56__rcx n1217__vss n164__i18__net5 n254__r_out n640__vss g45n2svt L=150e-9 W=6e-6 AD=1.2e-12 AS=1.2e-12 PD=12.4e-6 PS=12.4e-6 NRD=468.75e-3 NRS=468.75e-3 M=1
mi18__m15_55__rcx n319__r_out n218__i18__net5 n1191__vss n640__vss g45n2svt L=150e-9 W=6e-6 AD=1.2e-12 AS=1.2e-12 PD=12.4e-6 PS=12.4e-6 NRD=468.75e-3 NRS=468.75e-3 M=1
mi18__m15_54__rcx n1196__vss n214__i18__net5 n319__r_out n640__vss g45n2svt L=150e-9 W=6e-6 AD=1.2e-12 AS=1.2e-12 PD=12.4e-6 PS=12.4e-6 NRD=468.75e-3 NRS=468.75e-3 M=1
mi18__m15_53__rcx n306__r_out n208__i18__net5 n1196__vss n640__vss g45n2svt L=150e-9 W=6e-6 AD=1.2e-12 AS=1.2e-12 PD=12.4e-6 PS=12.4e-6 NRD=468.75e-3 NRS=468.75e-3 M=1
mi18__m15_52__rcx n1200__vss n203__i18__net5 n306__r_out n640__vss g45n2svt L=150e-9 W=6e-6 AD=1.2e-12 AS=1.2e-12 PD=12.4e-6 PS=12.4e-6 NRD=468.75e-3 NRS=468.75e-3 M=1
mi18__m15_51__rcx n293__r_out n199__i18__net5 n1200__vss n640__vss g45n2svt L=150e-9 W=6e-6 AD=1.2e-12 AS=1.2e-12 PD=12.4e-6 PS=12.4e-6 NRD=468.75e-3 NRS=468.75e-3 M=1
mi18__m15_50__rcx n1204__vss n193__i18__net5 n293__r_out n640__vss g45n2svt L=150e-9 W=6e-6 AD=1.2e-12 AS=1.2e-12 PD=12.4e-6 PS=12.4e-6 NRD=468.75e-3 NRS=468.75e-3 M=1
mi18__m15_49__rcx n356__r_out n250__i18__net5 n1179__vss n640__vss g45n2svt L=150e-9 W=6e-6 AD=1.2e-12 AS=1.2e-12 PD=12.4e-6 PS=12.4e-6 NRD=468.75e-3 NRS=468.75e-3 M=1
mi18__m15_48__rcx n1183__vss n245__i18__net5 n356__r_out n640__vss g45n2svt L=150e-9 W=6e-6 AD=1.2e-12 AS=1.2e-12 PD=12.4e-6 PS=12.4e-6 NRD=468.75e-3 NRS=468.75e-3 M=1
mi18__m15_47__rcx n339__r_out n240__i18__net5 n1183__vss n640__vss g45n2svt L=150e-9 W=6e-6 AD=1.2e-12 AS=1.2e-12 PD=12.4e-6 PS=12.4e-6 NRD=468.75e-3 NRS=468.75e-3 M=1
mi18__m15_46__rcx n1187__vss n235__i18__net5 n339__r_out n640__vss g45n2svt L=150e-9 W=6e-6 AD=1.2e-12 AS=1.2e-12 PD=12.4e-6 PS=12.4e-6 NRD=468.75e-3 NRS=468.75e-3 M=1
mi18__m15_45__rcx n332__r_out n228__i18__net5 n1187__vss n640__vss g45n2svt L=150e-9 W=6e-6 AD=1.2e-12 AS=1.2e-12 PD=12.4e-6 PS=12.4e-6 NRD=468.75e-3 NRS=468.75e-3 M=1
mi18__m15_44__rcx n1191__vss n223__i18__net5 n332__r_out n640__vss g45n2svt L=150e-9 W=6e-6 AD=1.2e-12 AS=1.2e-12 PD=12.4e-6 PS=12.4e-6 NRD=468.75e-3 NRS=468.75e-3 M=1
mi18__m15_43__rcx n395__r_out n278__i18__net5 n1167__vss n640__vss g45n2svt L=150e-9 W=6e-6 AD=1.2e-12 AS=1.2e-12 PD=12.4e-6 PS=12.4e-6 NRD=468.75e-3 NRS=468.75e-3 M=1
mi18__m15_42__rcx n1171__vss n275__i18__net5 n395__r_out n640__vss g45n2svt L=150e-9 W=6e-6 AD=1.2e-12 AS=1.2e-12 PD=12.4e-6 PS=12.4e-6 NRD=468.75e-3 NRS=468.75e-3 M=1
mi18__m15_41__rcx n382__r_out n268__i18__net5 n1171__vss n640__vss g45n2svt L=150e-9 W=6e-6 AD=1.2e-12 AS=1.2e-12 PD=12.4e-6 PS=12.4e-6 NRD=468.75e-3 NRS=468.75e-3 M=1
mi18__m15_40__rcx n1175__vss n265__i18__net5 n382__r_out n640__vss g45n2svt L=150e-9 W=6e-6 AD=1.2e-12 AS=1.2e-12 PD=12.4e-6 PS=12.4e-6 NRD=468.75e-3 NRS=468.75e-3 M=1
mi18__m15_39__rcx n371__r_out n258__i18__net5 n1175__vss n640__vss g45n2svt L=150e-9 W=6e-6 AD=1.2e-12 AS=1.2e-12 PD=12.4e-6 PS=12.4e-6 NRD=468.75e-3 NRS=468.75e-3 M=1
mi18__m15_38__rcx n1179__vss n253__i18__net5 n371__r_out n640__vss g45n2svt L=150e-9 W=6e-6 AD=1.2e-12 AS=1.2e-12 PD=12.4e-6 PS=12.4e-6 NRD=468.75e-3 NRS=468.75e-3 M=1
mi18__m15_37__rcx n1167__vss n283__i18__net5 n404__r_out n640__vss g45n2svt L=150e-9 W=6e-6 AD=1.2e-12 AS=1.2e-12 PD=12.4e-6 PS=12.4e-6 NRD=468.75e-3 NRS=468.75e-3 M=1
mi18__m15_36__rcx n1154__vss n313__i18__net5 n445__r_out n640__vss g45n2svt L=150e-9 W=6e-6 AD=1.2e-12 AS=1.2e-12 PD=12.4e-6 PS=12.4e-6 NRD=468.75e-3 NRS=468.75e-3 M=1
mi18__m15_35__rcx n438__r_out n310__i18__net5 n1154__vss n640__vss g45n2svt L=150e-9 W=6e-6 AD=1.2e-12 AS=1.2e-12 PD=12.4e-6 PS=12.4e-6 NRD=468.75e-3 NRS=468.75e-3 M=1
mi18__m15_34__rcx n1158__vss n303__i18__net5 n438__r_out n640__vss g45n2svt L=150e-9 W=6e-6 AD=1.2e-12 AS=1.2e-12 PD=12.4e-6 PS=12.4e-6 NRD=468.75e-3 NRS=468.75e-3 M=1
mi18__m15_33__rcx n417__r_out n298__i18__net5 n1158__vss n640__vss g45n2svt L=150e-9 W=6e-6 AD=1.2e-12 AS=1.2e-12 PD=12.4e-6 PS=12.4e-6 NRD=468.75e-3 NRS=468.75e-3 M=1
mi18__m15_32__rcx n1162__vss n293__i18__net5 n417__r_out n640__vss g45n2svt L=150e-9 W=6e-6 AD=1.2e-12 AS=1.2e-12 PD=12.4e-6 PS=12.4e-6 NRD=468.75e-3 NRS=468.75e-3 M=1
mi18__m15_31__rcx n404__r_out n288__i18__net5 n1162__vss n640__vss g45n2svt L=150e-9 W=6e-6 AD=1.2e-12 AS=1.2e-12 PD=12.4e-6 PS=12.4e-6 NRD=468.75e-3 NRS=468.75e-3 M=1
mi18__m15_30__rcx n1142__vss n345__i18__net5 n493__r_out n640__vss g45n2svt L=150e-9 W=6e-6 AD=1.2e-12 AS=1.2e-12 PD=12.4e-6 PS=12.4e-6 NRD=468.75e-3 NRS=468.75e-3 M=1
mi18__m15_29__rcx n478__r_out n338__i18__net5 n1142__vss n640__vss g45n2svt L=150e-9 W=6e-6 AD=1.2e-12 AS=1.2e-12 PD=12.4e-6 PS=12.4e-6 NRD=468.75e-3 NRS=468.75e-3 M=1
mi18__m15_28__rcx n1146__vss n335__i18__net5 n478__r_out n640__vss g45n2svt L=150e-9 W=6e-6 AD=1.2e-12 AS=1.2e-12 PD=12.4e-6 PS=12.4e-6 NRD=468.75e-3 NRS=468.75e-3 M=1
mi18__m15_27__rcx n461__r_out n328__i18__net5 n1146__vss n640__vss g45n2svt L=150e-9 W=6e-6 AD=1.2e-12 AS=1.2e-12 PD=12.4e-6 PS=12.4e-6 NRD=468.75e-3 NRS=468.75e-3 M=1
mi18__m15_26__rcx n1150__vss n325__i18__net5 n461__r_out n640__vss g45n2svt L=150e-9 W=6e-6 AD=1.2e-12 AS=1.2e-12 PD=12.4e-6 PS=12.4e-6 NRD=468.75e-3 NRS=468.75e-3 M=1
mi18__m15_25__rcx n445__r_out n320__i18__net5 n1150__vss n640__vss g45n2svt L=150e-9 W=6e-6 AD=1.2e-12 AS=1.2e-12 PD=12.4e-6 PS=12.4e-6 NRD=468.75e-3 NRS=468.75e-3 M=1
mi18__m15_24__rcx n1125__vss n375__i18__net5 n526__r_out n640__vss g45n2svt L=150e-9 W=6e-6 AD=1.2e-12 AS=1.2e-12 PD=12.4e-6 PS=12.4e-6 NRD=468.75e-3 NRS=468.75e-3 M=1
mi18__m15_23__rcx n517__r_out n368__i18__net5 n1125__vss n640__vss g45n2svt L=150e-9 W=6e-6 AD=1.2e-12 AS=1.2e-12 PD=12.4e-6 PS=12.4e-6 NRD=468.75e-3 NRS=468.75e-3 M=1
mi18__m15_22__rcx n1132__vss n365__i18__net5 n517__r_out n640__vss g45n2svt L=150e-9 W=6e-6 AD=1.2e-12 AS=1.2e-12 PD=12.4e-6 PS=12.4e-6 NRD=468.75e-3 NRS=468.75e-3 M=1
mi18__m15_21__rcx n506__r_out n360__i18__net5 n1132__vss n640__vss g45n2svt L=150e-9 W=6e-6 AD=1.2e-12 AS=1.2e-12 PD=12.4e-6 PS=12.4e-6 NRD=468.75e-3 NRS=468.75e-3 M=1
mi18__m15_20__rcx n1138__vss n355__i18__net5 n506__r_out n640__vss g45n2svt L=150e-9 W=6e-6 AD=1.2e-12 AS=1.2e-12 PD=12.4e-6 PS=12.4e-6 NRD=468.75e-3 NRS=468.75e-3 M=1
mi18__m15_19__rcx n493__r_out n348__i18__net5 n1138__vss n640__vss g45n2svt L=150e-9 W=6e-6 AD=1.2e-12 AS=1.2e-12 PD=12.4e-6 PS=12.4e-6 NRD=468.75e-3 NRS=468.75e-3 M=1
mi18__m15_18__rcx n1106__vss n405__i18__net5 n565__r_out n640__vss g45n2svt L=150e-9 W=6e-6 AD=1.2e-12 AS=1.2e-12 PD=12.4e-6 PS=12.4e-6 NRD=468.75e-3 NRS=468.75e-3 M=1
mi18__m15_17__rcx n552__r_out n398__i18__net5 n1106__vss n640__vss g45n2svt L=150e-9 W=6e-6 AD=1.2e-12 AS=1.2e-12 PD=12.4e-6 PS=12.4e-6 NRD=468.75e-3 NRS=468.75e-3 M=1
mi18__m15_16__rcx n1112__vss n395__i18__net5 n552__r_out n640__vss g45n2svt L=150e-9 W=6e-6 AD=1.2e-12 AS=1.2e-12 PD=12.4e-6 PS=12.4e-6 NRD=468.75e-3 NRS=468.75e-3 M=1
mi18__m15_15__rcx n539__r_out n390__i18__net5 n1112__vss n640__vss g45n2svt L=150e-9 W=6e-6 AD=1.2e-12 AS=1.2e-12 PD=12.4e-6 PS=12.4e-6 NRD=468.75e-3 NRS=468.75e-3 M=1
mi18__m15_14__rcx n1118__vss n385__i18__net5 n539__r_out n640__vss g45n2svt L=150e-9 W=6e-6 AD=1.2e-12 AS=1.2e-12 PD=12.4e-6 PS=12.4e-6 NRD=468.75e-3 NRS=468.75e-3 M=1
mi18__m15_13__rcx n526__r_out n378__i18__net5 n1118__vss n640__vss g45n2svt L=150e-9 W=6e-6 AD=1.2e-12 AS=1.2e-12 PD=12.4e-6 PS=12.4e-6 NRD=468.75e-3 NRS=468.75e-3 M=1
mi18__m15_12__rcx n565__r_out n408__i18__net5 n1098__vss n640__vss g45n2svt L=150e-9 W=6e-6 AD=1.2e-12 AS=1.2e-12 PD=12.4e-6 PS=12.4e-6 NRD=468.75e-3 NRS=468.75e-3 M=1
mi18__m15_11__rcx n604__r_out n440__i18__net5 n1081__vss n640__vss g45n2svt L=150e-9 W=6e-6 AD=1.2e-12 AS=1.2e-12 PD=12.4e-6 PS=12.4e-6 NRD=468.75e-3 NRS=468.75e-3 M=1
mi18__m15_10__rcx n1086__vss n435__i18__net5 n604__r_out n640__vss g45n2svt L=150e-9 W=6e-6 AD=1.2e-12 AS=1.2e-12 PD=12.4e-6 PS=12.4e-6 NRD=468.75e-3 NRS=468.75e-3 M=1
mi18__m15_9__rcx n591__r_out n428__i18__net5 n1086__vss n640__vss g45n2svt L=150e-9 W=6e-6 AD=1.2e-12 AS=1.2e-12 PD=12.4e-6 PS=12.4e-6 NRD=468.75e-3 NRS=468.75e-3 M=1
mi18__m15_8__rcx n1091__vss n423__i18__net5 n591__r_out n640__vss g45n2svt L=150e-9 W=6e-6 AD=1.2e-12 AS=1.2e-12 PD=12.4e-6 PS=12.4e-6 NRD=468.75e-3 NRS=468.75e-3 M=1
mi18__m15_7__rcx n578__r_out n419__i18__net5 n1091__vss n640__vss g45n2svt L=150e-9 W=6e-6 AD=1.2e-12 AS=1.2e-12 PD=12.4e-6 PS=12.4e-6 NRD=468.75e-3 NRS=468.75e-3 M=1
mi18__m15_6__rcx n1098__vss n413__i18__net5 n578__r_out n640__vss g45n2svt L=150e-9 W=6e-6 AD=1.2e-12 AS=1.2e-12 PD=12.4e-6 PS=12.4e-6 NRD=468.75e-3 NRS=468.75e-3 M=1
mi18__m15_5__rcx n1067__vss n463__i18__net5 n643__r_out n640__vss g45n2svt L=150e-9 W=6e-6 AD=1.2e-12 AS=1.2e-12 PD=12.4e-6 PS=12.4e-6 NRD=468.75e-3 NRS=468.75e-3 M=1
mi18__m15_4__rcx n630__r_out n458__i18__net5 n1067__vss n640__vss g45n2svt L=150e-9 W=6e-6 AD=1.2e-12 AS=1.2e-12 PD=12.4e-6 PS=12.4e-6 NRD=468.75e-3 NRS=468.75e-3 M=1
mi18__m15_3__rcx n1074__vss n453__i18__net5 n630__r_out n640__vss g45n2svt L=150e-9 W=6e-6 AD=1.2e-12 AS=1.2e-12 PD=12.4e-6 PS=12.4e-6 NRD=468.75e-3 NRS=468.75e-3 M=1
mi18__m15_2__rcx n617__r_out n450__i18__net5 n1074__vss n640__vss g45n2svt L=150e-9 W=6e-6 AD=1.2e-12 AS=1.2e-12 PD=12.4e-6 PS=12.4e-6 NRD=468.75e-3 NRS=468.75e-3 M=1
mi18__m15_1__rcx n1081__vss n443__i18__net5 n617__r_out n640__vss g45n2svt L=150e-9 W=6e-6 AD=1.2e-12 AS=1.2e-12 PD=12.4e-6 PS=12.4e-6 NRD=468.75e-3 NRS=468.75e-3 M=1
mi18__m15 n643__r_out n470__i18__net5 n1055__vss n640__vss g45n2svt L=150e-9 W=6e-6 AD=1.2e-12 AS=1.2e-12 PD=12.35e-6 PS=12.35e-6 NRD=468.75e-3 NRS=468.75e-3 M=1
mi18__m14_29__rcx n591__vss n19__i18__net4 n541__i18__net5 n640__vss g45n2svt L=150e-9 W=5.55e-6 AD=1.11e-12 AS=1.11e-12 PD=11.5e-6 PS=11.5e-6 NRD=468.75e-3 NRS=468.75e-3 M=1
mi18__m14_28__rcx n528__i18__net5 n16__i18__net4 n591__vss n640__vss g45n2svt L=150e-9 W=5.55e-6 AD=1.11e-12 AS=1.11e-12 PD=11.5e-6 PS=11.5e-6 NRD=468.75e-3 NRS=468.75e-3 M=1
mi18__m14_27__rcx n595__vss n13__i18__net4 n528__i18__net5 n640__vss g45n2svt L=150e-9 W=5.55e-6 AD=1.11e-12 AS=1.11e-12 PD=11.5e-6 PS=11.5e-6 NRD=468.75e-3 NRS=468.75e-3 M=1
mi18__m14_26__rcx n515__i18__net5 n10__i18__net4 n595__vss n640__vss g45n2svt L=150e-9 W=5.55e-6 AD=1.11e-12 AS=1.11e-12 PD=11.5e-6 PS=11.5e-6 NRD=468.75e-3 NRS=468.75e-3 M=1
mi18__m14_25__rcx n600__vss n7__i18__net4 n515__i18__net5 n640__vss g45n2svt L=150e-9 W=5.55e-6 AD=1.11e-12 AS=1.11e-12 PD=11.5e-6 PS=11.5e-6 NRD=468.75e-3 NRS=468.75e-3 M=1
mi18__m14_24__rcx n506__i18__net5 n4__i18__net4 n600__vss n640__vss g45n2svt L=150e-9 W=5.55e-6 AD=1.11e-12 AS=1.11e-12 PD=11.5e-6 PS=11.5e-6 NRD=468.75e-3 NRS=468.75e-3 M=1
mi18__m14_23__rcx n603__vss i18__net4 n506__i18__net5 n640__vss g45n2svt L=150e-9 W=5.55e-6 AD=832.5e-15 AS=832.5e-15 PD=11.45e-6 PS=11.45e-6 NRD=468.75e-3 NRS=468.75e-3 M=1
mi18__m14_22__rcx n580__i18__net5 n40__i18__net4 n572__vss n640__vss g45n2svt L=150e-9 W=5.55e-6 AD=1.11e-12 AS=1.11e-12 PD=11.5e-6 PS=11.5e-6 NRD=468.75e-3 NRS=468.75e-3 M=1
mi18__m14_21__rcx n577__vss n37__i18__net4 n580__i18__net5 n640__vss g45n2svt L=150e-9 W=5.55e-6 AD=1.11e-12 AS=1.11e-12 PD=11.5e-6 PS=11.5e-6 NRD=468.75e-3 NRS=468.75e-3 M=1
mi18__m14_20__rcx n567__i18__net5 n34__i18__net4 n577__vss n640__vss g45n2svt L=150e-9 W=5.55e-6 AD=1.11e-12 AS=1.11e-12 PD=11.5e-6 PS=11.5e-6 NRD=468.75e-3 NRS=468.75e-3 M=1
mi18__m14_19__rcx n583__vss n31__i18__net4 n567__i18__net5 n640__vss g45n2svt L=150e-9 W=5.55e-6 AD=1.11e-12 AS=1.11e-12 PD=11.5e-6 PS=11.5e-6 NRD=468.75e-3 NRS=468.75e-3 M=1
mi18__m14_18__rcx n560__i18__net5 n28__i18__net4 n583__vss n640__vss g45n2svt L=150e-9 W=5.55e-6 AD=1.11e-12 AS=1.11e-12 PD=11.5e-6 PS=11.5e-6 NRD=468.75e-3 NRS=468.75e-3 M=1
mi18__m14_17__rcx n587__vss n25__i18__net4 n560__i18__net5 n640__vss g45n2svt L=150e-9 W=5.55e-6 AD=1.11e-12 AS=1.11e-12 PD=11.5e-6 PS=11.5e-6 NRD=468.75e-3 NRS=468.75e-3 M=1
mi18__m14_16__rcx n541__i18__net5 n22__i18__net4 n587__vss n640__vss g45n2svt L=150e-9 W=5.55e-6 AD=1.11e-12 AS=1.11e-12 PD=11.5e-6 PS=11.5e-6 NRD=468.75e-3 NRS=468.75e-3 M=1
mi18__m14_15__rcx n572__vss n45__i18__net4 n599__i18__net5 n640__vss g45n2svt L=150e-9 W=5.55e-6 AD=1.11e-12 AS=1.11e-12 PD=11.5e-6 PS=11.5e-6 NRD=468.75e-3 NRS=468.75e-3 M=1
mi18__m14_14__rcx n638__i18__net5 n80__i18__net4 n555__vss n640__vss g45n2svt L=150e-9 W=5.55e-6 AD=1.11e-12 AS=1.11e-12 PD=11.5e-6 PS=11.5e-6 NRD=468.75e-3 NRS=468.75e-3 M=1
mi18__m14_13__rcx n559__vss n73__i18__net4 n638__i18__net5 n640__vss g45n2svt L=150e-9 W=5.55e-6 AD=1.11e-12 AS=1.11e-12 PD=11.5e-6 PS=11.5e-6 NRD=468.75e-3 NRS=468.75e-3 M=1
mi18__m14_12__rcx n619__i18__net5 n68__i18__net4 n559__vss n640__vss g45n2svt L=150e-9 W=5.55e-6 AD=1.11e-12 AS=1.11e-12 PD=11.5e-6 PS=11.5e-6 NRD=468.75e-3 NRS=468.75e-3 M=1
mi18__m14_11__rcx n564__vss n63__i18__net4 n619__i18__net5 n640__vss g45n2svt L=150e-9 W=5.55e-6 AD=1.11e-12 AS=1.11e-12 PD=11.5e-6 PS=11.5e-6 NRD=468.75e-3 NRS=468.75e-3 M=1
mi18__m14_10__rcx n606__i18__net5 n59__i18__net4 n564__vss n640__vss g45n2svt L=150e-9 W=5.55e-6 AD=1.11e-12 AS=1.11e-12 PD=11.5e-6 PS=11.5e-6 NRD=468.75e-3 NRS=468.75e-3 M=1
mi18__m14_9__rcx n568__vss n53__i18__net4 n606__i18__net5 n640__vss g45n2svt L=150e-9 W=5.55e-6 AD=1.11e-12 AS=1.11e-12 PD=11.5e-6 PS=11.5e-6 NRD=468.75e-3 NRS=468.75e-3 M=1
mi18__m14_8__rcx n599__i18__net5 n48__i18__net4 n568__vss n640__vss g45n2svt L=150e-9 W=5.55e-6 AD=1.11e-12 AS=1.11e-12 PD=11.5e-6 PS=11.5e-6 NRD=468.75e-3 NRS=468.75e-3 M=1
mi18__m14_7__rcx n542__vss n113__i18__net4 n684__i18__net5 n640__vss g45n2svt L=150e-9 W=5.55e-6 AD=1.11e-12 AS=1.11e-12 PD=11.5e-6 PS=11.5e-6 NRD=468.75e-3 NRS=468.75e-3 M=1
mi18__m14_6__rcx n677__i18__net5 n110__i18__net4 n542__vss n640__vss g45n2svt L=150e-9 W=5.55e-6 AD=1.11e-12 AS=1.11e-12 PD=11.5e-6 PS=11.5e-6 NRD=468.75e-3 NRS=468.75e-3 M=1
mi18__m14_5__rcx n547__vss n103__i18__net4 n677__i18__net5 n640__vss g45n2svt L=150e-9 W=5.55e-6 AD=1.11e-12 AS=1.11e-12 PD=11.5e-6 PS=11.5e-6 NRD=468.75e-3 NRS=468.75e-3 M=1
mi18__m14_4__rcx n658__i18__net5 n100__i18__net4 n547__vss n640__vss g45n2svt L=150e-9 W=5.55e-6 AD=1.11e-12 AS=1.11e-12 PD=11.5e-6 PS=11.5e-6 NRD=468.75e-3 NRS=468.75e-3 M=1
mi18__m14_3__rcx n551__vss n95__i18__net4 n658__i18__net5 n640__vss g45n2svt L=150e-9 W=5.55e-6 AD=1.11e-12 AS=1.11e-12 PD=11.5e-6 PS=11.5e-6 NRD=468.75e-3 NRS=468.75e-3 M=1
mi18__m14_2__rcx n645__i18__net5 n88__i18__net4 n551__vss n640__vss g45n2svt L=150e-9 W=5.55e-6 AD=1.11e-12 AS=1.11e-12 PD=11.5e-6 PS=11.5e-6 NRD=468.75e-3 NRS=468.75e-3 M=1
mi18__m14_1__rcx n555__vss n83__i18__net4 n645__i18__net5 n640__vss g45n2svt L=150e-9 W=5.55e-6 AD=1.11e-12 AS=1.11e-12 PD=11.5e-6 PS=11.5e-6 NRD=468.75e-3 NRS=468.75e-3 M=1
mi18__m3_9__rcx n196__i18__net4 n28__i18__net3 n623__vss n640__vss g45n2svt L=150e-9 W=4.58e-6 AD=916e-15 AS=916e-15 PD=9.51e-6 PS=9.51e-6 NRD=468.75e-3 NRS=468.75e-3 M=1
mi18__m3_8__rcx n629__vss n25__i18__net3 n196__i18__net4 n640__vss g45n2svt L=150e-9 W=4.58e-6 AD=916e-15 AS=916e-15 PD=9.56e-6 PS=9.56e-6 NRD=468.75e-3 NRS=468.75e-3 M=1
mi18__m3_7__rcx n185__i18__net4 n22__i18__net3 n629__vss n640__vss g45n2svt L=150e-9 W=4.58e-6 AD=916e-15 AS=916e-15 PD=9.56e-6 PS=9.56e-6 NRD=468.75e-3 NRS=468.75e-3 M=1
mi18__m3_6__rcx n631__vss n19__i18__net3 n185__i18__net4 n640__vss g45n2svt L=150e-9 W=4.58e-6 AD=916e-15 AS=916e-15 PD=9.56e-6 PS=9.56e-6 NRD=468.75e-3 NRS=468.75e-3 M=1
mi18__m3_5__rcx n180__i18__net4 n16__i18__net3 n631__vss n640__vss g45n2svt L=150e-9 W=4.58e-6 AD=916e-15 AS=916e-15 PD=9.56e-6 PS=9.56e-6 NRD=468.75e-3 NRS=468.75e-3 M=1
mi18__m3_4__rcx n633__vss n13__i18__net3 n180__i18__net4 n640__vss g45n2svt L=150e-9 W=4.58e-6 AD=916e-15 AS=916e-15 PD=9.56e-6 PS=9.56e-6 NRD=468.75e-3 NRS=468.75e-3 M=1
mi18__m3_3__rcx n163__i18__net4 n10__i18__net3 n633__vss n640__vss g45n2svt L=150e-9 W=4.58e-6 AD=916e-15 AS=916e-15 PD=9.56e-6 PS=9.56e-6 NRD=468.75e-3 NRS=468.75e-3 M=1
mi18__m3_2__rcx n636__vss n7__i18__net3 n163__i18__net4 n640__vss g45n2svt L=150e-9 W=4.58e-6 AD=916e-15 AS=916e-15 PD=9.56e-6 PS=9.56e-6 NRD=468.75e-3 NRS=468.75e-3 M=1
mi18__m3_1__rcx n152__i18__net4 n4__i18__net3 n636__vss n640__vss g45n2svt L=150e-9 W=4.58e-6 AD=916e-15 AS=916e-15 PD=9.56e-6 PS=9.56e-6 NRD=468.75e-3 NRS=468.75e-3 M=1
mi18__m3 n638__vss i18__net3 n152__i18__net4 n640__vss g45n2svt L=150e-9 W=4.58e-6 AD=687e-15 AS=687e-15 PD=9.51e-6 PS=9.51e-6 NRD=468.75e-3 NRS=468.75e-3 M=1
mi18__m14 n684__i18__net5 n120__i18__net4 n535__vss n640__vss g45n2svt L=150e-9 W=5.55e-6 AD=1.11e-12 AS=1.11e-12 PD=11.45e-6 PS=11.45e-6 NRD=468.75e-3 NRS=468.75e-3 M=1
mi18__m0 n7__i18__net1 serial_out_b_high_buff n1001__vss n640__vss g45n2svt L=150e-9 W=960e-9 AD=144e-15 AS=144e-15 PD=2.22e-6 PS=2.22e-6 NRD=468.75e-3 NRS=468.75e-3 M=1
mi18__m1_1__rcx n13__i18__net2 i18__net1 n1005__vss n640__vss g45n2svt L=150e-9 W=1.74e-6 AD=348e-15 AS=348e-15 PD=3.83e-6 PS=3.83e-6 NRD=468.75e-3 NRS=468.75e-3 M=1
mi18__m1 n1004__vss n6__i18__net1 n13__i18__net2 n640__vss g45n2svt L=150e-9 W=1.74e-6 AD=261e-15 AS=261e-15 PD=3.83e-6 PS=3.83e-6 NRD=468.75e-3 NRS=468.75e-3 M=1
mi18__m2_3__rcx n51__i18__net3 i18__net2 n708__vss n640__vss g45n2svt L=150e-9 W=3.16e-6 AD=632e-15 AS=632e-15 PD=6.67e-6 PS=6.67e-6 NRD=468.75e-3 NRS=468.75e-3 M=1
mi18__m2_2__rcx n711__vss n9__i18__net2 n51__i18__net3 n640__vss g45n2svt L=150e-9 W=3.16e-6 AD=632e-15 AS=632e-15 PD=6.72e-6 PS=6.72e-6 NRD=468.75e-3 NRS=468.75e-3 M=1
mi18__m2_1__rcx n60__i18__net3 n11__i18__net2 n711__vss n640__vss g45n2svt L=150e-9 W=3.16e-6 AD=632e-15 AS=632e-15 PD=6.72e-6 PS=6.72e-6 NRD=468.75e-3 NRS=468.75e-3 M=1
mi18__m2 n713__vss n12__i18__net2 n60__i18__net3 n640__vss g45n2svt L=150e-9 W=3.16e-6 AD=474e-15 AS=474e-15 PD=6.67e-6 PS=6.67e-6 NRD=468.75e-3 NRS=468.75e-3 M=1
mi12__nm0_2__rcx n9__i12__bio n6__i12__bcore_bar n1018__vss n640__vss g45n2svt L=150e-9 W=320e-9 AD=64e-15 AS=64e-15 PD=989.999e-9 PS=989.999e-9 NRD=468.75e-3 NRS=468.75e-3 M=1
mi12__nm0_1__rcx n1019__vss n4__i12__bcore_bar n9__i12__bio n640__vss g45n2svt L=150e-9 W=320e-9 AD=64e-15 AS=64e-15 PD=1.04e-6 PS=1.04e-6 NRD=468.75e-3 NRS=468.75e-3 M=1
mi12__nm0 n3__i12__bio n2__i12__bcore_bar n1019__vss n640__vss g45n2svt L=150e-9 W=320e-9 AD=48e-15 AS=48e-15 PD=989.999e-9 PS=989.999e-9 NRD=468.75e-3 NRS=468.75e-3 M=1
mi12__nm1_2__rcx n8__serial_out_b_high n6__serial_out n1021__vss n640__vss g45n2svt L=150e-9 W=320e-9 AD=64e-15 AS=64e-15 PD=989.999e-9 PS=989.999e-9 NRD=468.75e-3 NRS=468.75e-3 M=1
mi12__nm1_1__rcx n1023__vss n4__serial_out n8__serial_out_b_high n640__vss g45n2svt L=150e-9 W=320e-9 AD=64e-15 AS=64e-15 PD=1.04e-6 PS=1.04e-6 NRD=468.75e-3 NRS=468.75e-3 M=1
mi12__nm1 n10__serial_out_b_high n2__serial_out n1023__vss n640__vss g45n2svt L=150e-9 W=320e-9 AD=48e-15 AS=48e-15 PD=989.999e-9 PS=989.999e-9 NRD=468.75e-3 NRS=468.75e-3 M=1
mi36__m0_2__rcx n13__ck_buff n10__net13 n663__vss n640__vss g45n1svt L=45e-9 W=240e-9 AD=38.4e-15 AS=38.4e-15 PD=780e-9 PS=780e-9 NRD=1.16667 NRS=1.16667 M=1
mi36__m0_1__rcx n662__vss n8__net13 n13__ck_buff n640__vss g45n1svt L=45e-9 W=240e-9 AD=38.4e-15 AS=38.4e-15 PD=800e-9 PS=800e-9 NRD=1.16667 NRS=1.16667 M=1
mi36__m0 n24__ck_buff net13 n662__vss n640__vss g45n1svt L=45e-9 W=240e-9 AD=33.6e-15 AS=33.6e-15 PD=780e-9 PS=780e-9 NRD=1.16667 NRS=1.16667 M=1
mi32__m0_2__rcx n9__ck_b n6__net11 n668__vss n640__vss g45n1svt L=45e-9 W=240e-9 AD=38.4e-15 AS=38.4e-15 PD=780e-9 PS=780e-9 NRD=1.16667 NRS=1.16667 M=1
mi32__m0_1__rcx n669__vss n8__net11 n9__ck_b n640__vss g45n1svt L=45e-9 W=240e-9 AD=38.4e-15 AS=38.4e-15 PD=800e-9 PS=800e-9 NRD=1.16667 NRS=1.16667 M=1
mi32__m0 n5__ck_b n10__net11 n669__vss n640__vss g45n1svt L=45e-9 W=240e-9 AD=33.6e-15 AS=33.6e-15 PD=780e-9 PS=780e-9 NRD=1.16667 NRS=1.16667 M=1
mi37__m0_2__rcx n10__reset_buff n10__net14 n767__vss n640__vss g45n1svt L=45e-9 W=240e-9 AD=38.4e-15 AS=38.4e-15 PD=780e-9 PS=780e-9 NRD=1.16667 NRS=1.16667 M=1
mi37__m0_1__rcx n762__vss n8__net14 n10__reset_buff n640__vss g45n1svt L=45e-9 W=240e-9 AD=38.4e-15 AS=38.4e-15 PD=800e-9 PS=800e-9 NRD=1.16667 NRS=1.16667 M=1
mi37__m0 n13__reset_buff net14 n762__vss n640__vss g45n1svt L=45e-9 W=240e-9 AD=33.6e-15 AS=33.6e-15 PD=780e-9 PS=780e-9 NRD=1.16667 NRS=1.16667 M=1
mi33__m0_2__rcx n10__reset_b n6__net12 n790__vss n640__vss g45n1svt L=45e-9 W=240e-9 AD=38.4e-15 AS=38.4e-15 PD=780e-9 PS=780e-9 NRD=1.16667 NRS=1.16667 M=1
mi33__m0_1__rcx n793__vss n8__net12 n10__reset_b n640__vss g45n1svt L=45e-9 W=240e-9 AD=38.4e-15 AS=38.4e-15 PD=800e-9 PS=800e-9 NRD=1.16667 NRS=1.16667 M=1
mi33__m0 n7__reset_b n10__net12 n793__vss n640__vss g45n1svt L=45e-9 W=240e-9 AD=33.6e-15 AS=33.6e-15 PD=780e-9 PS=780e-9 NRD=1.16667 NRS=1.16667 M=1
mi30__m0_2__rcx n13__net11 n7__net9 n666__vss n640__vss g45n1svt L=45e-9 W=120e-9 AD=19.2e-15 AS=19.2e-15 PD=540e-9 PS=540e-9 NRD=1.16667 NRS=1.16667 M=1
mi30__m0_1__rcx n667__vss n9__net9 n13__net11 n640__vss g45n1svt L=45e-9 W=120e-9 AD=19.2e-15 AS=19.2e-15 PD=560e-9 PS=560e-9 NRD=1.16667 NRS=1.16667 M=1
mi30__m0 n18__net11 n10__net9 n667__vss n640__vss g45n1svt L=45e-9 W=120e-9 AD=16.8e-15 AS=16.8e-15 PD=540e-9 PS=540e-9 NRD=1.16667 NRS=1.16667 M=1
mi29__m0_2__rcx n15__r2_buff n10__net6 n733__vss n640__vss g45n1svt L=45e-9 W=120e-9 AD=19.2e-15 AS=19.2e-15 PD=540e-9 PS=540e-9 NRD=1.16667 NRS=1.16667 M=1
mi29__m0_1__rcx n732__vss n8__net6 n15__r2_buff n640__vss g45n1svt L=45e-9 W=120e-9 AD=19.2e-15 AS=19.2e-15 PD=560e-9 PS=560e-9 NRD=1.16667 NRS=1.16667 M=1
mi29__m0 n11__r2_buff net6 n732__vss n640__vss g45n1svt L=45e-9 W=120e-9 AD=16.8e-15 AS=16.8e-15 PD=540e-9 PS=540e-9 NRD=1.16667 NRS=1.16667 M=1
mi31__m0_2__rcx n13__net12 n7__net10 n782__vss n640__vss g45n1svt L=45e-9 W=120e-9 AD=19.2e-15 AS=19.2e-15 PD=540e-9 PS=540e-9 NRD=1.16667 NRS=1.16667 M=1
mi31__m0_1__rcx n787__vss n9__net10 n13__net12 n640__vss g45n1svt L=45e-9 W=120e-9 AD=19.2e-15 AS=19.2e-15 PD=560e-9 PS=560e-9 NRD=1.16667 NRS=1.16667 M=1
mi31__m0 n18__net12 n10__net10 n787__vss n640__vss g45n1svt L=45e-9 W=120e-9 AD=16.8e-15 AS=16.8e-15 PD=540e-9 PS=540e-9 NRD=1.16667 NRS=1.16667 M=1
mi27__m0_2__rcx n11__r0_buff n9__net7 n734__vss n640__vss g45n1svt L=45e-9 W=120e-9 AD=19.2e-15 AS=19.2e-15 PD=540e-9 PS=540e-9 NRD=1.16667 NRS=1.16667 M=1
mi27__m0_1__rcx n715__vss n7__net7 n11__r0_buff n640__vss g45n1svt L=45e-9 W=120e-9 AD=19.2e-15 AS=19.2e-15 PD=560e-9 PS=560e-9 NRD=1.16667 NRS=1.16667 M=1
mi27__m0 n13__r0_buff n6__net7 n715__vss n640__vss g45n1svt L=45e-9 W=120e-9 AD=16.8e-15 AS=16.8e-15 PD=540e-9 PS=540e-9 NRD=1.16667 NRS=1.16667 M=1
mi28__m0_2__rcx n11__r1_buff n9__net8 n941__vss n640__vss g45n1svt L=45e-9 W=120e-9 AD=19.2e-15 AS=19.2e-15 PD=540e-9 PS=540e-9 NRD=1.16667 NRS=1.16667 M=1
mi28__m0_1__rcx n887__vss n7__net8 n11__r1_buff n640__vss g45n1svt L=45e-9 W=120e-9 AD=19.2e-15 AS=19.2e-15 PD=560e-9 PS=560e-9 NRD=1.16667 NRS=1.16667 M=1
mi28__m0 n13__r1_buff n6__net8 n887__vss n640__vss g45n1svt L=45e-9 W=120e-9 AD=16.8e-15 AS=16.8e-15 PD=540e-9 PS=540e-9 NRD=1.16667 NRS=1.16667 M=1
mi34__m0 n14__net13 n26__ck n664__vss n640__vss g45n1svt L=45e-9 W=120e-9 AD=16.8e-15 AS=16.8e-15 PD=520e-9 PS=520e-9 NRD=1.16667 NRS=1.16667 M=1
mi16__m0 n11__net9 n25__ck n665__vss n640__vss g45n1svt L=45e-9 W=120e-9 AD=16.8e-15 AS=16.8e-15 PD=520e-9 PS=520e-9 NRD=1.16667 NRS=1.16667 M=1
mi23__m0 n13__net6 n5__r2 n735__vss n640__vss g45n1svt L=45e-9 W=120e-9 AD=16.8e-15 AS=16.8e-15 PD=520e-9 PS=520e-9 NRD=1.16667 NRS=1.16667 M=1
mi17__m0 n11__net10 n54__reset n776__vss n640__vss g45n1svt L=45e-9 W=120e-9 AD=16.8e-15 AS=16.8e-15 PD=520e-9 PS=520e-9 NRD=1.16667 NRS=1.16667 M=1
mi35__m0 n11__net14 n55__reset n771__vss n640__vss g45n1svt L=45e-9 W=120e-9 AD=16.8e-15 AS=16.8e-15 PD=520e-9 PS=520e-9 NRD=1.16667 NRS=1.16667 M=1
mi19__m0 n12__net7 n13__r0 n736__vss n640__vss g45n1svt L=45e-9 W=120e-9 AD=16.8e-15 AS=16.8e-15 PD=520e-9 PS=520e-9 NRD=1.16667 NRS=1.16667 M=1
mi22__m0 n12__net8 n4__r1 n942__vss n640__vss g45n1svt L=45e-9 W=120e-9 AD=16.8e-15 AS=16.8e-15 PD=520e-9 PS=520e-9 NRD=1.16667 NRS=1.16667 M=1
mi2__nm18 n752__vss n21__reset_buff n14__i2__net74 n640__vss g45n1svt L=45e-9 W=120e-9 AD=16.8e-15 AS=16.8e-15 PD=520e-9 PS=520e-9 NRD=1.16667 NRS=1.16667 M=1
mi2__nm2_1__rcx n9__i2__net75 n6__i2__net74 n750__vss n640__vss g45n1svt L=45e-9 W=240e-9 AD=38.4e-15 AS=38.4e-15 PD=780e-9 PS=780e-9 NRD=1.16667 NRS=1.16667 M=1
mi2__nm2 n748__vss n5__i2__net74 n9__i2__net75 n640__vss g45n1svt L=45e-9 W=240e-9 AD=33.6e-15 AS=33.6e-15 PD=780e-9 PS=780e-9 NRD=1.16667 NRS=1.16667 M=1
mi2__nm12 n12__i2__net76 n29__ck_buff n10__i2__net75 n640__vss g45n1svt L=45e-9 W=120e-9 AD=16.8e-15 AS=16.8e-15 PD=520e-9 PS=520e-9 NRD=1.16667 NRS=1.16667 M=1
mi2__nm15 n746__vss n2__i2__net77 n8__i2__net76 n640__vss g45n1svt L=570e-9 W=120e-9 AD=16.8e-15 AS=16.8e-15 PD=520e-9 PS=520e-9 NRD=1.16667 NRS=1.16667 M=1
mi2__nm13_1__rcx n8__i2__net77 n6__i2__net76 n744__vss n640__vss g45n1svt L=45e-9 W=240e-9 AD=38.4e-15 AS=38.4e-15 PD=780e-9 PS=780e-9 NRD=1.16667 NRS=1.16667 M=1
mi2__nm13 n742__vss n5__i2__net76 n8__i2__net77 n640__vss g45n1svt L=45e-9 W=240e-9 AD=33.6e-15 AS=33.6e-15 PD=780e-9 PS=780e-9 NRD=1.16667 NRS=1.16667 M=1
mi2__nm16 n21__serial_out n6__i2__net77 n740__vss n640__vss g45n1svt L=45e-9 W=240e-9 AD=33.6e-15 AS=33.6e-15 PD=760e-9 PS=760e-9 NRD=1.16667 NRS=1.16667 M=1
mi2__nm17 n3__i2__q n10__serial_out n738__vss n640__vss g45n1svt L=45e-9 W=240e-9 AD=33.6e-15 AS=33.6e-15 PD=760e-9 PS=760e-9 NRD=1.16667 NRS=1.16667 M=1
mi2__nm21 n6__i2__net79 n4__shift n763__vss n640__vss g45n1svt L=45e-9 W=120e-9 AD=16.8e-15 AS=16.8e-15 PD=520e-9 PS=520e-9 NRD=1.16667 NRS=1.16667 M=1
mi2__nm22 n7__i2__net1 n13__shift n5__net4 n640__vss g45n1svt L=45e-9 W=120e-9 AD=19.2e-15 AS=19.2e-15 PD=540e-9 PS=540e-9 NRD=1.16667 NRS=1.16667 M=1
mi2__nm20 n5__r0_buff n3__i2__net79 n7__i2__net1 n640__vss g45n1svt L=45e-9 W=120e-9 AD=16.8e-15 AS=16.8e-15 PD=540e-9 PS=540e-9 NRD=1.16667 NRS=1.16667 M=1
mi2__nm1 n4__i2__net73 n4__i2__net1 n759__vss n640__vss g45n1svt L=45e-9 W=240e-9 AD=33.6e-15 AS=33.6e-15 PD=760e-9 PS=760e-9 NRD=1.16667 NRS=1.16667 M=1
mi2__nm0 n12__i2__net74 n20__ck_b n5__i2__net73 n640__vss g45n1svt L=45e-9 W=120e-9 AD=16.8e-15 AS=16.8e-15 PD=520e-9 PS=520e-9 NRD=1.16667 NRS=1.16667 M=1
mi2__nm8 n756__vss n2__i2__net75 n8__i2__net74 n640__vss g45n1svt L=570e-9 W=120e-9 AD=16.8e-15 AS=16.8e-15 PD=520e-9 PS=520e-9 NRD=1.16667 NRS=1.16667 M=1
mi1__nm18 n751__vss n23__reset_buff n14__i1__net74 n640__vss g45n1svt L=45e-9 W=120e-9 AD=16.8e-15 AS=16.8e-15 PD=520e-9 PS=520e-9 NRD=1.16667 NRS=1.16667 M=1
mi1__nm2_1__rcx n12__i1__net75 n7__i1__net74 n749__vss n640__vss g45n1svt L=45e-9 W=240e-9 AD=38.4e-15 AS=38.4e-15 PD=780e-9 PS=780e-9 NRD=1.16667 NRS=1.16667 M=1
mi1__nm2 n747__vss i1__net74 n12__i1__net75 n640__vss g45n1svt L=45e-9 W=240e-9 AD=33.6e-15 AS=33.6e-15 PD=780e-9 PS=780e-9 NRD=1.16667 NRS=1.16667 M=1
mi1__nm12 n13__i1__net76 n31__ck_buff n6__i1__net75 n640__vss g45n1svt L=45e-9 W=120e-9 AD=16.8e-15 AS=16.8e-15 PD=520e-9 PS=520e-9 NRD=1.16667 NRS=1.16667 M=1
mi1__nm15 n745__vss n3__i1__net77 n8__i1__net76 n640__vss g45n1svt L=570e-9 W=120e-9 AD=16.8e-15 AS=16.8e-15 PD=520e-9 PS=520e-9 NRD=1.16667 NRS=1.16667 M=1
mi1__nm13_1__rcx n8__i1__net77 n7__i1__net76 n743__vss n640__vss g45n1svt L=45e-9 W=240e-9 AD=38.4e-15 AS=38.4e-15 PD=780e-9 PS=780e-9 NRD=1.16667 NRS=1.16667 M=1
mi1__nm13 n741__vss i1__net76 n8__i1__net77 n640__vss g45n1svt L=45e-9 W=240e-9 AD=33.6e-15 AS=33.6e-15 PD=780e-9 PS=780e-9 NRD=1.16667 NRS=1.16667 M=1
mi1__nm16 n15__net4 n4__i1__net77 n739__vss n640__vss g45n1svt L=45e-9 W=240e-9 AD=33.6e-15 AS=33.6e-15 PD=760e-9 PS=760e-9 NRD=1.16667 NRS=1.16667 M=1
mi1__nm17 i1__q n8__net4 n737__vss n640__vss g45n1svt L=45e-9 W=240e-9 AD=33.6e-15 AS=33.6e-15 PD=760e-9 PS=760e-9 NRD=1.16667 NRS=1.16667 M=1
mi1__nm21 n6__i1__net79 n5__shift n758__vss n640__vss g45n1svt L=45e-9 W=120e-9 AD=16.8e-15 AS=16.8e-15 PD=520e-9 PS=520e-9 NRD=1.16667 NRS=1.16667 M=1
mi1__nm22 n7__i1__net1 n15__shift n5__net3 n640__vss g45n1svt L=45e-9 W=120e-9 AD=19.2e-15 AS=19.2e-15 PD=540e-9 PS=540e-9 NRD=1.16667 NRS=1.16667 M=1
mi1__nm20 n5__r1_buff n3__i1__net79 n7__i1__net1 n640__vss g45n1svt L=45e-9 W=120e-9 AD=16.8e-15 AS=16.8e-15 PD=540e-9 PS=540e-9 NRD=1.16667 NRS=1.16667 M=1
mi1__nm1 n6__i1__net73 i1__net1 n755__vss n640__vss g45n1svt L=45e-9 W=240e-9 AD=33.6e-15 AS=33.6e-15 PD=760e-9 PS=760e-9 NRD=1.16667 NRS=1.16667 M=1
mi1__nm0 n13__i1__net74 n22__ck_b i1__net73 n640__vss g45n1svt L=45e-9 W=120e-9 AD=16.8e-15 AS=16.8e-15 PD=520e-9 PS=520e-9 NRD=1.16667 NRS=1.16667 M=1
mi1__nm8 n753__vss n3__i1__net75 n8__i1__net74 n640__vss g45n1svt L=570e-9 W=120e-9 AD=16.8e-15 AS=16.8e-15 PD=520e-9 PS=520e-9 NRD=1.16667 NRS=1.16667 M=1
mi0__nm18 n952__vss n25__reset_buff n14__i0__net74 n640__vss g45n1svt L=45e-9 W=120e-9 AD=16.8e-15 AS=16.8e-15 PD=520e-9 PS=520e-9 NRD=1.16667 NRS=1.16667 M=1
mi0__nm2_1__rcx n9__i0__net75 n6__i0__net74 n950__vss n640__vss g45n1svt L=45e-9 W=240e-9 AD=38.4e-15 AS=38.4e-15 PD=780e-9 PS=780e-9 NRD=1.16667 NRS=1.16667 M=1
mi0__nm2 n948__vss n5__i0__net74 n9__i0__net75 n640__vss g45n1svt L=45e-9 W=240e-9 AD=33.6e-15 AS=33.6e-15 PD=780e-9 PS=780e-9 NRD=1.16667 NRS=1.16667 M=1
mi0__nm12 n12__i0__net76 n33__ck_buff n10__i0__net75 n640__vss g45n1svt L=45e-9 W=120e-9 AD=16.8e-15 AS=16.8e-15 PD=520e-9 PS=520e-9 NRD=1.16667 NRS=1.16667 M=1
mi0__nm15 n947__vss n2__i0__net77 n8__i0__net76 n640__vss g45n1svt L=570e-9 W=120e-9 AD=16.8e-15 AS=16.8e-15 PD=520e-9 PS=520e-9 NRD=1.16667 NRS=1.16667 M=1
mi0__nm13_1__rcx n8__i0__net77 n6__i0__net76 n946__vss n640__vss g45n1svt L=45e-9 W=240e-9 AD=38.4e-15 AS=38.4e-15 PD=780e-9 PS=780e-9 NRD=1.16667 NRS=1.16667 M=1
mi0__nm13 n945__vss n5__i0__net76 n8__i0__net77 n640__vss g45n1svt L=45e-9 W=240e-9 AD=33.6e-15 AS=33.6e-15 PD=780e-9 PS=780e-9 NRD=1.16667 NRS=1.16667 M=1
mi0__nm16 n11__net3 n6__i0__net77 n944__vss n640__vss g45n1svt L=45e-9 W=240e-9 AD=33.6e-15 AS=33.6e-15 PD=760e-9 PS=760e-9 NRD=1.16667 NRS=1.16667 M=1
mi0__nm17 n3__i0__q n9__net3 n943__vss n640__vss g45n1svt L=45e-9 W=240e-9 AD=33.6e-15 AS=33.6e-15 PD=760e-9 PS=760e-9 NRD=1.16667 NRS=1.16667 M=1
mi0__nm21 n6__i0__net79 n12__shift n959__vss n640__vss g45n1svt L=45e-9 W=120e-9 AD=16.8e-15 AS=16.8e-15 PD=520e-9 PS=520e-9 NRD=1.16667 NRS=1.16667 M=1
mi0__nm22 n7__i0__net1 n17__shift n529__vss n640__vss g45n1svt L=45e-9 W=120e-9 AD=19.2e-15 AS=19.2e-15 PD=540e-9 PS=540e-9 NRD=1.16667 NRS=1.16667 M=1
mi0__nm20 n5__r2_buff n3__i0__net79 n7__i0__net1 n640__vss g45n1svt L=45e-9 W=120e-9 AD=16.8e-15 AS=16.8e-15 PD=540e-9 PS=540e-9 NRD=1.16667 NRS=1.16667 M=1
mi0__nm1 n4__i0__net73 n4__i0__net1 n955__vss n640__vss g45n1svt L=45e-9 W=240e-9 AD=33.6e-15 AS=33.6e-15 PD=760e-9 PS=760e-9 NRD=1.16667 NRS=1.16667 M=1
mi0__nm0 n12__i0__net74 n24__ck_b n5__i0__net73 n640__vss g45n1svt L=45e-9 W=120e-9 AD=16.8e-15 AS=16.8e-15 PD=520e-9 PS=520e-9 NRD=1.16667 NRS=1.16667 M=1
mi0__nm8 n953__vss n2__i0__net75 n8__i0__net74 n640__vss g45n1svt L=570e-9 W=120e-9 AD=16.8e-15 AS=16.8e-15 PD=520e-9 PS=520e-9 NRD=1.16667 NRS=1.16667 M=1
mi14__nm0_5__rcx n672__vss n23__i14__net7 n86__i14__net9 n640__vss g45n1svt L=45e-9 W=240e-9 AD=38.4e-15 AS=38.4e-15 PD=800e-9 PS=800e-9 NRD=1.16667 NRS=1.16667 M=1
mi14__nm0_4__rcx n89__i14__net9 n21__i14__net7 n672__vss n640__vss g45n1svt L=45e-9 W=240e-9 AD=38.4e-15 AS=38.4e-15 PD=800e-9 PS=800e-9 NRD=1.16667 NRS=1.16667 M=1
mi14__nm0_3__rcx n671__vss n19__i14__net7 n89__i14__net9 n640__vss g45n1svt L=45e-9 W=240e-9 AD=38.4e-15 AS=38.4e-15 PD=800e-9 PS=800e-9 NRD=1.16667 NRS=1.16667 M=1
mi14__nm0_2__rcx n92__i14__net9 n17__i14__net7 n671__vss n640__vss g45n1svt L=45e-9 W=240e-9 AD=38.4e-15 AS=38.4e-15 PD=800e-9 PS=800e-9 NRD=1.16667 NRS=1.16667 M=1
mi14__nm0_1__rcx n670__vss n5__i14__net7 n92__i14__net9 n640__vss g45n1svt L=45e-9 W=240e-9 AD=33.6e-15 AS=33.6e-15 PD=780e-9 PS=780e-9 NRD=1.16667 NRS=1.16667 M=1
mi14__nm0 n86__i14__net9 n24__i14__net7 n673__vss n640__vss g45n1svt L=45e-9 W=240e-9 AD=38.4e-15 AS=38.4e-15 PD=780e-9 PS=780e-9 NRD=1.16667 NRS=1.16667 M=1
mi14__nm8_5__rcx n679__vss n44__reset n49__i14__net4 n640__vss g45n1svt L=45e-9 W=240e-9 AD=38.4e-15 AS=38.4e-15 PD=800e-9 PS=800e-9 NRD=1.16667 NRS=1.16667 M=1
mi14__nm8_4__rcx n52__i14__net4 n42__reset n679__vss n640__vss g45n1svt L=45e-9 W=240e-9 AD=38.4e-15 AS=38.4e-15 PD=800e-9 PS=800e-9 NRD=1.16667 NRS=1.16667 M=1
mi14__nm8_3__rcx n678__vss n40__reset n52__i14__net4 n640__vss g45n1svt L=45e-9 W=240e-9 AD=38.4e-15 AS=38.4e-15 PD=800e-9 PS=800e-9 NRD=1.16667 NRS=1.16667 M=1
mi14__nm8_2__rcx n55__i14__net4 n38__reset n678__vss n640__vss g45n1svt L=45e-9 W=240e-9 AD=38.4e-15 AS=38.4e-15 PD=800e-9 PS=800e-9 NRD=1.16667 NRS=1.16667 M=1
mi14__nm8_1__rcx n676__vss n26__reset n55__i14__net4 n640__vss g45n1svt L=45e-9 W=240e-9 AD=33.6e-15 AS=33.6e-15 PD=780e-9 PS=780e-9 NRD=1.16667 NRS=1.16667 M=1
mi14__nm8 n49__i14__net4 n45__reset n681__vss n640__vss g45n1svt L=45e-9 W=240e-9 AD=38.4e-15 AS=38.4e-15 PD=780e-9 PS=780e-9 NRD=1.16667 NRS=1.16667 M=1
mi14__nm1_5__rcx n814__vss n22__i14__net11 n99__i14__net10 n640__vss g45n1svt L=45e-9 W=240e-9 AD=38.4e-15 AS=38.4e-15 PD=800e-9 PS=800e-9 NRD=1.16667 NRS=1.16667 M=1
mi14__nm1_4__rcx n102__i14__net10 n20__i14__net11 n814__vss n640__vss g45n1svt L=45e-9 W=240e-9 AD=38.4e-15 AS=38.4e-15 PD=800e-9 PS=800e-9 NRD=1.16667 NRS=1.16667 M=1
mi14__nm1_3__rcx n810__vss n18__i14__net11 n102__i14__net10 n640__vss g45n1svt L=45e-9 W=240e-9 AD=38.4e-15 AS=38.4e-15 PD=800e-9 PS=800e-9 NRD=1.16667 NRS=1.16667 M=1
mi14__nm1_2__rcx n105__i14__net10 n16__i14__net11 n810__vss n640__vss g45n1svt L=45e-9 W=240e-9 AD=38.4e-15 AS=38.4e-15 PD=800e-9 PS=800e-9 NRD=1.16667 NRS=1.16667 M=1
mi14__nm1_1__rcx n806__vss n15__i14__net11 n105__i14__net10 n640__vss g45n1svt L=45e-9 W=240e-9 AD=33.6e-15 AS=33.6e-15 PD=780e-9 PS=780e-9 NRD=1.16667 NRS=1.16667 M=1
mi14__nm1 n99__i14__net10 n14__i14__net11 n818__vss n640__vss g45n1svt L=45e-9 W=240e-9 AD=38.4e-15 AS=38.4e-15 PD=780e-9 PS=780e-9 NRD=1.16667 NRS=1.16667 M=1
mi14__nm7_5__rcx n831__vss n46__i14__net4 n59__i14__net3 n640__vss g45n1svt L=45e-9 W=240e-9 AD=38.4e-15 AS=38.4e-15 PD=800e-9 PS=800e-9 NRD=1.16667 NRS=1.16667 M=1
mi14__nm7_4__rcx n62__i14__net3 n44__i14__net4 n831__vss n640__vss g45n1svt L=45e-9 W=240e-9 AD=38.4e-15 AS=38.4e-15 PD=800e-9 PS=800e-9 NRD=1.16667 NRS=1.16667 M=1
mi14__nm7_3__rcx n830__vss n42__i14__net4 n62__i14__net3 n640__vss g45n1svt L=45e-9 W=240e-9 AD=38.4e-15 AS=38.4e-15 PD=800e-9 PS=800e-9 NRD=1.16667 NRS=1.16667 M=1
mi14__nm7_2__rcx n71__i14__net3 n40__i14__net4 n830__vss n640__vss g45n1svt L=45e-9 W=240e-9 AD=38.4e-15 AS=38.4e-15 PD=800e-9 PS=800e-9 NRD=1.16667 NRS=1.16667 M=1
mi14__nm7_1__rcx n822__vss n39__i14__net4 n71__i14__net3 n640__vss g45n1svt L=45e-9 W=240e-9 AD=33.6e-15 AS=33.6e-15 PD=780e-9 PS=780e-9 NRD=1.16667 NRS=1.16667 M=1
mi14__nm7 n59__i14__net3 n38__i14__net4 n832__vss n640__vss g45n1svt L=45e-9 W=240e-9 AD=38.4e-15 AS=38.4e-15 PD=780e-9 PS=780e-9 NRD=1.16667 NRS=1.16667 M=1
mi14__i17__i2__nm0 n13__i14__i17__i2__net1 n2__i14__i17__net3 n5__i14__i17__net1 n640__vss g45n1svt L=45e-9 W=120e-9 AD=16.8e-15 AS=16.8e-15 PD=520e-9 PS=520e-9 NRD=1.16667 NRS=1.16667 M=1
mi14__i17__i2__nm8 n705__vss n3__i14__i17__i2__net2 n8__i14__i17__i2__net1 n640__vss g45n1svt L=570e-9 W=120e-9 AD=16.8e-15 AS=16.8e-15 PD=520e-9 PS=520e-9 NRD=1.16667 NRS=1.16667 M=1
mi14__i17__i2__nm18 n703__vss n5__reset n15__i14__i17__i2__net1 n640__vss g45n1svt L=45e-9 W=120e-9 AD=16.8e-15 AS=16.8e-15 PD=520e-9 PS=520e-9 NRD=1.16667 NRS=1.16667 M=1
mi14__i17__i2__nm2_1__rcx n12__i14__i17__i2__net2 n7__i14__i17__i2__net1 n701__vss n640__vss g45n1svt L=45e-9 W=240e-9 AD=38.4e-15 AS=38.4e-15 PD=780e-9 PS=780e-9 NRD=1.16667 NRS=1.16667 M=1
mi14__i17__i2__nm2 n699__vss i14__i17__i2__net1 n12__i14__i17__i2__net2 n640__vss g45n1svt L=45e-9 W=240e-9 AD=33.6e-15 AS=33.6e-15 PD=780e-9 PS=780e-9 NRD=1.16667 NRS=1.16667 M=1
mi14__i17__i2__nm12 n13__i14__i17__i2__net5 n7__ck n6__i14__i17__i2__net2 n640__vss g45n1svt L=45e-9 W=120e-9 AD=16.8e-15 AS=16.8e-15 PD=520e-9 PS=520e-9 NRD=1.16667 NRS=1.16667 M=1
mi14__i17__i2__nm15 n696__vss n3__i14__i17__i2__net4 n8__i14__i17__i2__net5 n640__vss g45n1svt L=570e-9 W=120e-9 AD=16.8e-15 AS=16.8e-15 PD=520e-9 PS=520e-9 NRD=1.16667 NRS=1.16667 M=1
mi14__i17__i2__nm13_1__rcx n8__i14__i17__i2__net4 n7__i14__i17__i2__net5 n694__vss n640__vss g45n1svt L=45e-9 W=240e-9 AD=38.4e-15 AS=38.4e-15 PD=780e-9 PS=780e-9 NRD=1.16667 NRS=1.16667 M=1
mi14__i17__i2__nm13 n692__vss i14__i17__i2__net5 n8__i14__i17__i2__net4 n640__vss g45n1svt L=45e-9 W=240e-9 AD=33.6e-15 AS=33.6e-15 PD=780e-9 PS=780e-9 NRD=1.16667 NRS=1.16667 M=1
mi14__i17__i2__nm16 n29__i14__i17__net1 n4__i14__i17__i2__net4 n690__vss n640__vss g45n1svt L=45e-9 W=240e-9 AD=33.6e-15 AS=33.6e-15 PD=760e-9 PS=760e-9 NRD=1.16667 NRS=1.16667 M=1
mi14__i17__i2__nm17 n17__i14__i17__net7 n14__i14__i17__net1 n688__vss n640__vss g45n1svt L=45e-9 W=240e-9 AD=33.6e-15 AS=33.6e-15 PD=760e-9 PS=760e-9 NRD=1.16667 NRS=1.16667 M=1
mi14__i17__i3__nm0 n12__i14__i17__i3__net1 n2__i14__i17__net1 n3__i14__i17__net8 n640__vss g45n1svt L=45e-9 W=120e-9 AD=16.8e-15 AS=16.8e-15 PD=520e-9 PS=520e-9 NRD=1.16667 NRS=1.16667 M=1
mi14__i17__i3__nm8 n885__vss n2__i14__i17__i3__net2 n8__i14__i17__i3__net1 n640__vss g45n1svt L=570e-9 W=120e-9 AD=16.8e-15 AS=16.8e-15 PD=520e-9 PS=520e-9 NRD=1.16667 NRS=1.16667 M=1
mi14__i17__i3__nm18 n880__vss n7__reset n15__i14__i17__i3__net1 n640__vss g45n1svt L=45e-9 W=120e-9 AD=16.8e-15 AS=16.8e-15 PD=520e-9 PS=520e-9 NRD=1.16667 NRS=1.16667 M=1
mi14__i17__i3__nm2_1__rcx n9__i14__i17__i3__net2 n6__i14__i17__i3__net1 n876__vss n640__vss g45n1svt L=45e-9 W=240e-9 AD=38.4e-15 AS=38.4e-15 PD=780e-9 PS=780e-9 NRD=1.16667 NRS=1.16667 M=1
mi14__i17__i3__nm2 n875__vss n5__i14__i17__i3__net1 n9__i14__i17__i3__net2 n640__vss g45n1svt L=45e-9 W=240e-9 AD=33.6e-15 AS=33.6e-15 PD=780e-9 PS=780e-9 NRD=1.16667 NRS=1.16667 M=1
mi14__i17__i3__nm12 n12__i14__i17__i3__net5 n4__i14__i17__net7 n10__i14__i17__i3__net2 n640__vss g45n1svt L=45e-9 W=120e-9 AD=16.8e-15 AS=16.8e-15 PD=520e-9 PS=520e-9 NRD=1.16667 NRS=1.16667 M=1
mi14__i17__i3__nm15 n867__vss n2__i14__i17__i3__net4 n8__i14__i17__i3__net5 n640__vss g45n1svt L=570e-9 W=120e-9 AD=16.8e-15 AS=16.8e-15 PD=520e-9 PS=520e-9 NRD=1.16667 NRS=1.16667 M=1
mi14__i17__i3__nm13_1__rcx n8__i14__i17__i3__net4 n6__i14__i17__i3__net5 n863__vss n640__vss g45n1svt L=45e-9 W=240e-9 AD=38.4e-15 AS=38.4e-15 PD=780e-9 PS=780e-9 NRD=1.16667 NRS=1.16667 M=1
mi14__i17__i3__nm13 n859__vss n5__i14__i17__i3__net5 n8__i14__i17__i3__net4 n640__vss g45n1svt L=45e-9 W=240e-9 AD=33.6e-15 AS=33.6e-15 PD=780e-9 PS=780e-9 NRD=1.16667 NRS=1.16667 M=1
mi14__i17__i3__nm16 n20__i14__i17__net8 n6__i14__i17__i3__net4 n858__vss n640__vss g45n1svt L=45e-9 W=240e-9 AD=33.6e-15 AS=33.6e-15 PD=760e-9 PS=760e-9 NRD=1.16667 NRS=1.16667 M=1
mi14__i17__i3__nm17 n12__i14__i17__net11 n9__i14__i17__net8 n854__vss n640__vss g45n1svt L=45e-9 W=240e-9 AD=33.6e-15 AS=33.6e-15 PD=760e-9 PS=760e-9 NRD=1.16667 NRS=1.16667 M=1
mi14__i17__i4__nm3 n10__i14__i17__net9 n3__i14__i17__net11 n851__vss n640__vss g45n1svt L=45e-9 W=120e-9 AD=19.2e-15 AS=19.2e-15 PD=540e-9 PS=540e-9 NRD=1.16667 NRS=1.16667 M=1
mi14__i17__i4__nm2 n270__vdd n13__i14__i17__net8 n10__i14__i17__net9 n640__vss g45n1svt L=45e-9 W=120e-9 AD=16.8e-15 AS=16.8e-15 PD=540e-9 PS=540e-9 NRD=1.16667 NRS=1.16667 M=1
mi14__i17__i4__nm6 n13__i14__i17__net10 n7__i14__i17__net9 n850__vss n640__vss g45n1svt L=45e-9 W=240e-9 AD=33.6e-15 AS=33.6e-15 PD=760e-9 PS=760e-9 NRD=1.16667 NRS=1.16667 M=1
mi14__i17__i4__nm5 n841__vss n7__i14__i17__net10 n20__i14__i17__net9 n640__vss g45n1svt L=45e-9 W=240e-9 AD=33.6e-15 AS=33.6e-15 PD=760e-9 PS=760e-9 NRD=1.16667 NRS=1.16667 M=1
mi14__i17__i4__nm1 n20__i14__i17__net10 n4__i14__i17__net11 n262__vdd n640__vss g45n1svt L=45e-9 W=120e-9 AD=19.2e-15 AS=19.2e-15 PD=540e-9 PS=540e-9 NRD=1.16667 NRS=1.16667 M=1
mi14__i17__i4__nm0 n833__vss n14__i14__i17__net8 n20__i14__i17__net10 n640__vss g45n1svt L=45e-9 W=120e-9 AD=16.8e-15 AS=16.8e-15 PD=540e-9 PS=540e-9 NRD=1.16667 NRS=1.16667 M=1
mi14__i17__nm0 n5__i14__i17__net3 n1__ck n707__vss n640__vss g45n1svt L=45e-9 W=120e-9 AD=16.8e-15 AS=16.8e-15 PD=520e-9 PS=520e-9 NRD=1.16667 NRS=1.16667 M=1
mi14__i17__nm1 n7__i14__i17__net6 n3__reset n886__vss n640__vss g45n1svt L=45e-9 W=120e-9 AD=16.8e-15 AS=16.8e-15 PD=520e-9 PS=520e-9 NRD=1.16667 NRS=1.16667 M=1
mi14__i17__nm14 n25__i14__net11 i14__i17__net10 n685__vss n640__vss g45n1svt L=45e-9 W=240e-9 AD=33.6e-15 AS=33.6e-15 PD=760e-9 PS=760e-9 NRD=1.16667 NRS=1.16667 M=1
mi14__i17__nm15 n26__i14__net7 i14__i17__net9 n683__vss n640__vss g45n1svt L=45e-9 W=240e-9 AD=33.6e-15 AS=33.6e-15 PD=760e-9 PS=760e-9 NRD=1.16667 NRS=1.16667 M=1
mi14__i11__nm0 n13__i14__i11__net1 n34__i14__net9 n1__y3 n640__vss g45n1svt L=45e-9 W=120e-9 AD=16.8e-15 AS=16.8e-15 PD=520e-9 PS=520e-9 NRD=1.16667 NRS=1.16667 M=1
mi14__i11__nm8 n843__vss n3__i14__i11__net2 n8__i14__i11__net1 n640__vss g45n1svt L=570e-9 W=120e-9 AD=16.8e-15 AS=16.8e-15 PD=520e-9 PS=520e-9 NRD=1.16667 NRS=1.16667 M=1
mi14__i11__nm18 n840__vss n30__i14__net3 n15__i14__i11__net1 n640__vss g45n1svt L=45e-9 W=120e-9 AD=16.8e-15 AS=16.8e-15 PD=520e-9 PS=520e-9 NRD=1.16667 NRS=1.16667 M=1
mi14__i11__nm2_1__rcx n12__i14__i11__net2 n7__i14__i11__net1 n836__vss n640__vss g45n1svt L=45e-9 W=240e-9 AD=38.4e-15 AS=38.4e-15 PD=780e-9 PS=780e-9 NRD=1.16667 NRS=1.16667 M=1
mi14__i11__nm2 n829__vss i14__i11__net1 n12__i14__i11__net2 n640__vss g45n1svt L=45e-9 W=240e-9 AD=33.6e-15 AS=33.6e-15 PD=780e-9 PS=780e-9 NRD=1.16667 NRS=1.16667 M=1
mi14__i11__nm12 n13__i14__i11__net5 n58__i14__net10 n6__i14__i11__net2 n640__vss g45n1svt L=45e-9 W=120e-9 AD=16.8e-15 AS=16.8e-15 PD=520e-9 PS=520e-9 NRD=1.16667 NRS=1.16667 M=1
mi14__i11__nm15 n821__vss n3__i14__i11__net4 n8__i14__i11__net5 n640__vss g45n1svt L=570e-9 W=120e-9 AD=16.8e-15 AS=16.8e-15 PD=520e-9 PS=520e-9 NRD=1.16667 NRS=1.16667 M=1
mi14__i11__nm13_1__rcx n9__i14__i11__net4 n7__i14__i11__net5 n817__vss n640__vss g45n1svt L=45e-9 W=240e-9 AD=38.4e-15 AS=38.4e-15 PD=780e-9 PS=780e-9 NRD=1.16667 NRS=1.16667 M=1
mi14__i11__nm13 n813__vss i14__i11__net5 n9__i14__i11__net4 n640__vss g45n1svt L=45e-9 W=240e-9 AD=33.6e-15 AS=33.6e-15 PD=780e-9 PS=780e-9 NRD=1.16667 NRS=1.16667 M=1
mi14__i11__nm16 n10__i14__x_out_b_1 n4__i14__i11__net4 n809__vss n640__vss g45n1svt L=45e-9 W=240e-9 AD=33.6e-15 AS=33.6e-15 PD=760e-9 PS=760e-9 NRD=1.16667 NRS=1.16667 M=1
mi14__i11__nm17 n7__y_out_3 i14__x_out_b_1 n801__vss n640__vss g45n1svt L=45e-9 W=240e-9 AD=33.6e-15 AS=33.6e-15 PD=760e-9 PS=760e-9 NRD=1.16667 NRS=1.16667 M=1
mi14__i13__nm0 n13__i14__i13__net1 n2__i14__net9 n1__x3 n640__vss g45n1svt L=45e-9 W=120e-9 AD=16.8e-15 AS=16.8e-15 PD=520e-9 PS=520e-9 NRD=1.16667 NRS=1.16667 M=1
mi14__i13__nm8 n884__vss n3__i14__i13__net2 n8__i14__i13__net1 n640__vss g45n1svt L=570e-9 W=120e-9 AD=16.8e-15 AS=16.8e-15 PD=520e-9 PS=520e-9 NRD=1.16667 NRS=1.16667 M=1
mi14__i13__nm18 n882__vss n2__i14__net3 n15__i14__i13__net1 n640__vss g45n1svt L=45e-9 W=120e-9 AD=16.8e-15 AS=16.8e-15 PD=520e-9 PS=520e-9 NRD=1.16667 NRS=1.16667 M=1
mi14__i13__nm2_1__rcx n12__i14__i13__net2 n7__i14__i13__net1 n879__vss n640__vss g45n1svt L=45e-9 W=240e-9 AD=38.4e-15 AS=38.4e-15 PD=780e-9 PS=780e-9 NRD=1.16667 NRS=1.16667 M=1
mi14__i13__nm2 n874__vss i14__i13__net1 n12__i14__i13__net2 n640__vss g45n1svt L=45e-9 W=240e-9 AD=33.6e-15 AS=33.6e-15 PD=780e-9 PS=780e-9 NRD=1.16667 NRS=1.16667 M=1
mi14__i13__nm12 n13__i14__i13__net5 n10__i14__net10 n6__i14__i13__net2 n640__vss g45n1svt L=45e-9 W=120e-9 AD=16.8e-15 AS=16.8e-15 PD=520e-9 PS=520e-9 NRD=1.16667 NRS=1.16667 M=1
mi14__i13__nm15 n869__vss n3__i14__i13__net4 n8__i14__i13__net5 n640__vss g45n1svt L=570e-9 W=120e-9 AD=16.8e-15 AS=16.8e-15 PD=520e-9 PS=520e-9 NRD=1.16667 NRS=1.16667 M=1
mi14__i13__nm13_1__rcx n8__i14__i13__net4 n7__i14__i13__net5 n866__vss n640__vss g45n1svt L=45e-9 W=240e-9 AD=38.4e-15 AS=38.4e-15 PD=780e-9 PS=780e-9 NRD=1.16667 NRS=1.16667 M=1
mi14__i13__nm13 n862__vss i14__i13__net5 n8__i14__i13__net4 n640__vss g45n1svt L=45e-9 W=240e-9 AD=33.6e-15 AS=33.6e-15 PD=780e-9 PS=780e-9 NRD=1.16667 NRS=1.16667 M=1
mi14__i13__nm16 n10__i14__y_out_b_3 n4__i14__i13__net4 n857__vss n640__vss g45n1svt L=45e-9 W=240e-9 AD=33.6e-15 AS=33.6e-15 PD=760e-9 PS=760e-9 NRD=1.16667 NRS=1.16667 M=1
mi14__i13__nm17 x_out_3 i14__y_out_b_3 n849__vss n640__vss g45n1svt L=45e-9 W=240e-9 AD=33.6e-15 AS=33.6e-15 PD=760e-9 PS=760e-9 NRD=1.16667 NRS=1.16667 M=1
mi14__i15__nm0 n13__i14__i15__net1 n38__i14__net9 n1__y1 n640__vss g45n1svt L=45e-9 W=120e-9 AD=16.8e-15 AS=16.8e-15 PD=520e-9 PS=520e-9 NRD=1.16667 NRS=1.16667 M=1
mi14__i15__nm8 n981__vss n3__i14__i15__net2 n8__i14__i15__net1 n640__vss g45n1svt L=570e-9 W=120e-9 AD=16.8e-15 AS=16.8e-15 PD=520e-9 PS=520e-9 NRD=1.16667 NRS=1.16667 M=1
mi14__i15__nm18 n979__vss n34__i14__net3 n15__i14__i15__net1 n640__vss g45n1svt L=45e-9 W=120e-9 AD=16.8e-15 AS=16.8e-15 PD=520e-9 PS=520e-9 NRD=1.16667 NRS=1.16667 M=1
mi14__i15__nm2_1__rcx n12__i14__i15__net2 n7__i14__i15__net1 n977__vss n640__vss g45n1svt L=45e-9 W=240e-9 AD=38.4e-15 AS=38.4e-15 PD=780e-9 PS=780e-9 NRD=1.16667 NRS=1.16667 M=1
mi14__i15__nm2 n975__vss i14__i15__net1 n12__i14__i15__net2 n640__vss g45n1svt L=45e-9 W=240e-9 AD=33.6e-15 AS=33.6e-15 PD=780e-9 PS=780e-9 NRD=1.16667 NRS=1.16667 M=1
mi14__i15__nm12 n13__i14__i15__net5 n62__i14__net10 n6__i14__i15__net2 n640__vss g45n1svt L=45e-9 W=120e-9 AD=16.8e-15 AS=16.8e-15 PD=520e-9 PS=520e-9 NRD=1.16667 NRS=1.16667 M=1
mi14__i15__nm15 n973__vss n3__i14__i15__net4 n8__i14__i15__net5 n640__vss g45n1svt L=570e-9 W=120e-9 AD=16.8e-15 AS=16.8e-15 PD=520e-9 PS=520e-9 NRD=1.16667 NRS=1.16667 M=1
mi14__i15__nm13_1__rcx n9__i14__i15__net4 n7__i14__i15__net5 n971__vss n640__vss g45n1svt L=45e-9 W=240e-9 AD=38.4e-15 AS=38.4e-15 PD=780e-9 PS=780e-9 NRD=1.16667 NRS=1.16667 M=1
mi14__i15__nm13 n969__vss i14__i15__net5 n9__i14__i15__net4 n640__vss g45n1svt L=45e-9 W=240e-9 AD=33.6e-15 AS=33.6e-15 PD=780e-9 PS=780e-9 NRD=1.16667 NRS=1.16667 M=1
mi14__i15__nm16 n10__i14__y_out_b_1 n4__i14__i15__net4 n967__vss n640__vss g45n1svt L=45e-9 W=240e-9 AD=33.6e-15 AS=33.6e-15 PD=760e-9 PS=760e-9 NRD=1.16667 NRS=1.16667 M=1
mi14__i15__nm17 n7__y_out_1 i14__y_out_b_1 n965__vss n640__vss g45n1svt L=45e-9 W=240e-9 AD=33.6e-15 AS=33.6e-15 PD=760e-9 PS=760e-9 NRD=1.16667 NRS=1.16667 M=1
mi14__i10__nm0 n13__i14__i10__net1 n6__i14__net9 n1__x1 n640__vss g45n1svt L=45e-9 W=120e-9 AD=16.8e-15 AS=16.8e-15 PD=520e-9 PS=520e-9 NRD=1.16667 NRS=1.16667 M=1
mi14__i10__nm8 n999__vss n3__i14__i10__net2 n8__i14__i10__net1 n640__vss g45n1svt L=570e-9 W=120e-9 AD=16.8e-15 AS=16.8e-15 PD=520e-9 PS=520e-9 NRD=1.16667 NRS=1.16667 M=1
mi14__i10__nm18 n997__vss n6__i14__net3 n15__i14__i10__net1 n640__vss g45n1svt L=45e-9 W=120e-9 AD=16.8e-15 AS=16.8e-15 PD=520e-9 PS=520e-9 NRD=1.16667 NRS=1.16667 M=1
mi14__i10__nm2_1__rcx n12__i14__i10__net2 n7__i14__i10__net1 n995__vss n640__vss g45n1svt L=45e-9 W=240e-9 AD=38.4e-15 AS=38.4e-15 PD=780e-9 PS=780e-9 NRD=1.16667 NRS=1.16667 M=1
mi14__i10__nm2 n993__vss i14__i10__net1 n12__i14__i10__net2 n640__vss g45n1svt L=45e-9 W=240e-9 AD=33.6e-15 AS=33.6e-15 PD=780e-9 PS=780e-9 NRD=1.16667 NRS=1.16667 M=1
mi14__i10__nm12 n13__i14__i10__net5 n14__i14__net10 n6__i14__i10__net2 n640__vss g45n1svt L=45e-9 W=120e-9 AD=16.8e-15 AS=16.8e-15 PD=520e-9 PS=520e-9 NRD=1.16667 NRS=1.16667 M=1
mi14__i10__nm15 n991__vss n3__i14__i10__net4 n8__i14__i10__net5 n640__vss g45n1svt L=570e-9 W=120e-9 AD=16.8e-15 AS=16.8e-15 PD=520e-9 PS=520e-9 NRD=1.16667 NRS=1.16667 M=1
mi14__i10__nm13_1__rcx n8__i14__i10__net4 n7__i14__i10__net5 n989__vss n640__vss g45n1svt L=45e-9 W=240e-9 AD=38.4e-15 AS=38.4e-15 PD=780e-9 PS=780e-9 NRD=1.16667 NRS=1.16667 M=1
mi14__i10__nm13 n987__vss i14__i10__net5 n8__i14__i10__net4 n640__vss g45n1svt L=45e-9 W=240e-9 AD=33.6e-15 AS=33.6e-15 PD=780e-9 PS=780e-9 NRD=1.16667 NRS=1.16667 M=1
mi14__i10__nm16 n10__i14__x_out_b_2 n4__i14__i10__net4 n985__vss n640__vss g45n1svt L=45e-9 W=240e-9 AD=33.6e-15 AS=33.6e-15 PD=760e-9 PS=760e-9 NRD=1.16667 NRS=1.16667 M=1
mi14__i10__nm17 x_out_1 i14__x_out_b_2 n983__vss n640__vss g45n1svt L=45e-9 W=240e-9 AD=33.6e-15 AS=33.6e-15 PD=760e-9 PS=760e-9 NRD=1.16667 NRS=1.16667 M=1
mi14__i14__nm0 n12__i14__i14__net1 n36__i14__net9 n3__y2 n640__vss g45n1svt L=45e-9 W=120e-9 AD=16.8e-15 AS=16.8e-15 PD=520e-9 PS=520e-9 NRD=1.16667 NRS=1.16667 M=1
mi14__i14__nm8 n982__vss n2__i14__i14__net2 n8__i14__i14__net1 n640__vss g45n1svt L=570e-9 W=120e-9 AD=16.8e-15 AS=16.8e-15 PD=520e-9 PS=520e-9 NRD=1.16667 NRS=1.16667 M=1
mi14__i14__nm18 n980__vss n32__i14__net3 n15__i14__i14__net1 n640__vss g45n1svt L=45e-9 W=120e-9 AD=16.8e-15 AS=16.8e-15 PD=520e-9 PS=520e-9 NRD=1.16667 NRS=1.16667 M=1
mi14__i14__nm2_1__rcx n9__i14__i14__net2 n6__i14__i14__net1 n978__vss n640__vss g45n1svt L=45e-9 W=240e-9 AD=38.4e-15 AS=38.4e-15 PD=780e-9 PS=780e-9 NRD=1.16667 NRS=1.16667 M=1
mi14__i14__nm2 n976__vss n5__i14__i14__net1 n9__i14__i14__net2 n640__vss g45n1svt L=45e-9 W=240e-9 AD=33.6e-15 AS=33.6e-15 PD=780e-9 PS=780e-9 NRD=1.16667 NRS=1.16667 M=1
mi14__i14__nm12 n12__i14__i14__net5 n60__i14__net10 n10__i14__i14__net2 n640__vss g45n1svt L=45e-9 W=120e-9 AD=16.8e-15 AS=16.8e-15 PD=520e-9 PS=520e-9 NRD=1.16667 NRS=1.16667 M=1
mi14__i14__nm15 n974__vss n2__i14__i14__net4 n8__i14__i14__net5 n640__vss g45n1svt L=570e-9 W=120e-9 AD=16.8e-15 AS=16.8e-15 PD=520e-9 PS=520e-9 NRD=1.16667 NRS=1.16667 M=1
mi14__i14__nm13_1__rcx n9__i14__i14__net4 n6__i14__i14__net5 n972__vss n640__vss g45n1svt L=45e-9 W=240e-9 AD=38.4e-15 AS=38.4e-15 PD=780e-9 PS=780e-9 NRD=1.16667 NRS=1.16667 M=1
mi14__i14__nm13 n970__vss n5__i14__i14__net5 n9__i14__i14__net4 n640__vss g45n1svt L=45e-9 W=240e-9 AD=33.6e-15 AS=33.6e-15 PD=780e-9 PS=780e-9 NRD=1.16667 NRS=1.16667 M=1
mi14__i14__nm16 n8__i14__y_out_b_2 n6__i14__i14__net4 n968__vss n640__vss g45n1svt L=45e-9 W=240e-9 AD=33.6e-15 AS=33.6e-15 PD=760e-9 PS=760e-9 NRD=1.16667 NRS=1.16667 M=1
mi14__i14__nm17 n9__y_out_2 n4__i14__y_out_b_2 n966__vss n640__vss g45n1svt L=45e-9 W=240e-9 AD=33.6e-15 AS=33.6e-15 PD=760e-9 PS=760e-9 NRD=1.16667 NRS=1.16667 M=1
mi14__i16__nm0 n12__i14__i16__net1 n4__i14__net9 n3__x2 n640__vss g45n1svt L=45e-9 W=120e-9 AD=16.8e-15 AS=16.8e-15 PD=520e-9 PS=520e-9 NRD=1.16667 NRS=1.16667 M=1
mi14__i16__nm8 n1000__vss n2__i14__i16__net2 n8__i14__i16__net1 n640__vss g45n1svt L=570e-9 W=120e-9 AD=16.8e-15 AS=16.8e-15 PD=520e-9 PS=520e-9 NRD=1.16667 NRS=1.16667 M=1
mi14__i16__nm18 n998__vss n4__i14__net3 n15__i14__i16__net1 n640__vss g45n1svt L=45e-9 W=120e-9 AD=16.8e-15 AS=16.8e-15 PD=520e-9 PS=520e-9 NRD=1.16667 NRS=1.16667 M=1
mi14__i16__nm2_1__rcx n9__i14__i16__net2 n6__i14__i16__net1 n996__vss n640__vss g45n1svt L=45e-9 W=240e-9 AD=38.4e-15 AS=38.4e-15 PD=780e-9 PS=780e-9 NRD=1.16667 NRS=1.16667 M=1
mi14__i16__nm2 n994__vss n5__i14__i16__net1 n9__i14__i16__net2 n640__vss g45n1svt L=45e-9 W=240e-9 AD=33.6e-15 AS=33.6e-15 PD=780e-9 PS=780e-9 NRD=1.16667 NRS=1.16667 M=1
mi14__i16__nm12 n12__i14__i16__net5 n12__i14__net10 n10__i14__i16__net2 n640__vss g45n1svt L=45e-9 W=120e-9 AD=16.8e-15 AS=16.8e-15 PD=520e-9 PS=520e-9 NRD=1.16667 NRS=1.16667 M=1
mi14__i16__nm15 n992__vss n2__i14__i16__net4 n8__i14__i16__net5 n640__vss g45n1svt L=570e-9 W=120e-9 AD=16.8e-15 AS=16.8e-15 PD=520e-9 PS=520e-9 NRD=1.16667 NRS=1.16667 M=1
mi14__i16__nm13_1__rcx n8__i14__i16__net4 n6__i14__i16__net5 n990__vss n640__vss g45n1svt L=45e-9 W=240e-9 AD=38.4e-15 AS=38.4e-15 PD=780e-9 PS=780e-9 NRD=1.16667 NRS=1.16667 M=1
mi14__i16__nm13 n988__vss n5__i14__i16__net5 n8__i14__i16__net4 n640__vss g45n1svt L=45e-9 W=240e-9 AD=33.6e-15 AS=33.6e-15 PD=780e-9 PS=780e-9 NRD=1.16667 NRS=1.16667 M=1
mi14__i16__nm16 n8__i14__y_out_b_0 n6__i14__i16__net4 n986__vss n640__vss g45n1svt L=45e-9 W=240e-9 AD=33.6e-15 AS=33.6e-15 PD=760e-9 PS=760e-9 NRD=1.16667 NRS=1.16667 M=1
mi14__i16__nm17 n3__x_out_2 n4__i14__y_out_b_0 n984__vss n640__vss g45n1svt L=45e-9 W=240e-9 AD=33.6e-15 AS=33.6e-15 PD=760e-9 PS=760e-9 NRD=1.16667 NRS=1.16667 M=1
mi14__i12__nm0 n12__i14__i12__net1 n40__i14__net9 n3__y0 n640__vss g45n1svt L=45e-9 W=120e-9 AD=16.8e-15 AS=16.8e-15 PD=520e-9 PS=520e-9 NRD=1.16667 NRS=1.16667 M=1
mi14__i12__nm8 n1084__vss n2__i14__i12__net2 n8__i14__i12__net1 n640__vss g45n1svt L=570e-9 W=120e-9 AD=16.8e-15 AS=16.8e-15 PD=520e-9 PS=520e-9 NRD=1.16667 NRS=1.16667 M=1
mi14__i12__nm18 n1078__vss n36__i14__net3 n15__i14__i12__net1 n640__vss g45n1svt L=45e-9 W=120e-9 AD=16.8e-15 AS=16.8e-15 PD=520e-9 PS=520e-9 NRD=1.16667 NRS=1.16667 M=1
mi14__i12__nm2_1__rcx n9__i14__i12__net2 n6__i14__i12__net1 n1077__vss n640__vss g45n1svt L=45e-9 W=240e-9 AD=38.4e-15 AS=38.4e-15 PD=780e-9 PS=780e-9 NRD=1.16667 NRS=1.16667 M=1
mi14__i12__nm2 n1070__vss n5__i14__i12__net1 n9__i14__i12__net2 n640__vss g45n1svt L=45e-9 W=240e-9 AD=33.6e-15 AS=33.6e-15 PD=780e-9 PS=780e-9 NRD=1.16667 NRS=1.16667 M=1
mi14__i12__nm12 n12__i14__i12__net5 n64__i14__net10 n10__i14__i12__net2 n640__vss g45n1svt L=45e-9 W=120e-9 AD=16.8e-15 AS=16.8e-15 PD=520e-9 PS=520e-9 NRD=1.16667 NRS=1.16667 M=1
mi14__i12__nm15 n1064__vss n2__i14__i12__net4 n8__i14__i12__net5 n640__vss g45n1svt L=570e-9 W=120e-9 AD=16.8e-15 AS=16.8e-15 PD=520e-9 PS=520e-9 NRD=1.16667 NRS=1.16667 M=1
mi14__i12__nm13_1__rcx n9__i14__i12__net4 n6__i14__i12__net5 n1063__vss n640__vss g45n1svt L=45e-9 W=240e-9 AD=38.4e-15 AS=38.4e-15 PD=780e-9 PS=780e-9 NRD=1.16667 NRS=1.16667 M=1
mi14__i12__nm13 n1062__vss n5__i14__i12__net5 n9__i14__i12__net4 n640__vss g45n1svt L=45e-9 W=240e-9 AD=33.6e-15 AS=33.6e-15 PD=780e-9 PS=780e-9 NRD=1.16667 NRS=1.16667 M=1
mi14__i12__nm16 n8__i14__x_out_b_0 n6__i14__i12__net4 n1061__vss n640__vss g45n1svt L=45e-9 W=240e-9 AD=33.6e-15 AS=33.6e-15 PD=760e-9 PS=760e-9 NRD=1.16667 NRS=1.16667 M=1
mi14__i12__nm17 n11__y_out_0 n4__i14__x_out_b_0 n1060__vss n640__vss g45n1svt L=45e-9 W=240e-9 AD=33.6e-15 AS=33.6e-15 PD=760e-9 PS=760e-9 NRD=1.16667 NRS=1.16667 M=1
mi14__i9__nm0 n12__i14__i9__net1 n8__i14__net9 n3__x0 n640__vss g45n1svt L=45e-9 W=120e-9 AD=16.8e-15 AS=16.8e-15 PD=520e-9 PS=520e-9 NRD=1.16667 NRS=1.16667 M=1
mi14__i9__nm8 n1135__vss n2__i14__i9__net2 n8__i14__i9__net1 n640__vss g45n1svt L=570e-9 W=120e-9 AD=16.8e-15 AS=16.8e-15 PD=520e-9 PS=520e-9 NRD=1.16667 NRS=1.16667 M=1
mi14__i9__nm18 n1129__vss n8__i14__net3 n15__i14__i9__net1 n640__vss g45n1svt L=45e-9 W=120e-9 AD=16.8e-15 AS=16.8e-15 PD=520e-9 PS=520e-9 NRD=1.16667 NRS=1.16667 M=1
mi14__i9__nm2_1__rcx n9__i14__i9__net2 n6__i14__i9__net1 n1128__vss n640__vss g45n1svt L=45e-9 W=240e-9 AD=38.4e-15 AS=38.4e-15 PD=780e-9 PS=780e-9 NRD=1.16667 NRS=1.16667 M=1
mi14__i9__nm2 n1121__vss n5__i14__i9__net1 n9__i14__i9__net2 n640__vss g45n1svt L=45e-9 W=240e-9 AD=33.6e-15 AS=33.6e-15 PD=780e-9 PS=780e-9 NRD=1.16667 NRS=1.16667 M=1
mi14__i9__nm12 n12__i14__i9__net5 n16__i14__net10 n10__i14__i9__net2 n640__vss g45n1svt L=45e-9 W=120e-9 AD=16.8e-15 AS=16.8e-15 PD=520e-9 PS=520e-9 NRD=1.16667 NRS=1.16667 M=1
mi14__i9__nm15 n1110__vss n2__i14__i9__net4 n8__i14__i9__net5 n640__vss g45n1svt L=570e-9 W=120e-9 AD=16.8e-15 AS=16.8e-15 PD=520e-9 PS=520e-9 NRD=1.16667 NRS=1.16667 M=1
mi14__i9__nm13_1__rcx n8__i14__i9__net4 n6__i14__i9__net5 n1109__vss n640__vss g45n1svt L=45e-9 W=240e-9 AD=38.4e-15 AS=38.4e-15 PD=780e-9 PS=780e-9 NRD=1.16667 NRS=1.16667 M=1
mi14__i9__nm13 n1102__vss n5__i14__i9__net5 n8__i14__i9__net4 n640__vss g45n1svt L=45e-9 W=240e-9 AD=33.6e-15 AS=33.6e-15 PD=780e-9 PS=780e-9 NRD=1.16667 NRS=1.16667 M=1
mi14__i9__nm16 n8__i14__x_out_b_3 n6__i14__i9__net4 n1101__vss n640__vss g45n1svt L=45e-9 W=240e-9 AD=33.6e-15 AS=33.6e-15 PD=760e-9 PS=760e-9 NRD=1.16667 NRS=1.16667 M=1
mi14__i9__nm17 n3__x_out_0 n4__i14__x_out_b_3 n1094__vss n640__vss g45n1svt L=45e-9 W=240e-9 AD=33.6e-15 AS=33.6e-15 PD=760e-9 PS=760e-9 NRD=1.16667 NRS=1.16667 M=1
mi14__nm10 n2__i14__clk_div4_out_b i14__net7 n675__vss n640__vss g45n1svt L=45e-9 W=240e-9 AD=33.6e-15 AS=33.6e-15 PD=760e-9 PS=760e-9 NRD=1.16667 NRS=1.16667 M=1
mi14__nm9 ck4 i14__net11 n674__vss n640__vss g45n1svt L=45e-9 W=240e-9 AD=33.6e-15 AS=33.6e-15 PD=760e-9 PS=760e-9 NRD=1.16667 NRS=1.16667 M=1
mi13__i20__i4__nm2 n3__i13__i20__i4__net2 n5__i13__net18 n949__vss n640__vss g45n1svt L=45e-9 W=120e-9 AD=16.8e-15 AS=16.8e-15 PD=520e-9 PS=520e-9 NRD=1.16667 NRS=1.16667 M=1
mi13__i20__i4__nm0 n5__r1 i13__i20__i4__net2 n16__i13__net7 n640__vss g45n1svt L=45e-9 W=120e-9 AD=16.8e-15 AS=16.8e-15 PD=520e-9 PS=520e-9 NRD=1.16667 NRS=1.16667 M=1
mi13__i20__i4__nm1 n9__r1 n5__i13__net7 n10__i13__i20__i4__net2 n640__vss g45n1svt L=45e-9 W=120e-9 AD=16.8e-15 AS=16.8e-15 PD=520e-9 PS=520e-9 NRD=1.16667 NRS=1.16667 M=1
mi13__i20__nm0 n8__i13__i20__net1 i13__net18 i13__i20__net3 n640__vss g45n1svt L=45e-9 W=240e-9 AD=33.6e-15 AS=33.6e-15 PD=780e-9 PS=780e-9 NRD=1.16667 NRS=1.16667 M=1
mi13__i20__nm1 i13__i20__net3 i13__net7 n954__vss n640__vss g45n1svt L=45e-9 W=240e-9 AD=38.4e-15 AS=38.4e-15 PD=780e-9 PS=780e-9 NRD=1.16667 NRS=1.16667 M=1
mi13__i20__nm3 n7__i13__net23 i13__i20__net1 n951__vss n640__vss g45n1svt L=45e-9 W=120e-9 AD=16.8e-15 AS=16.8e-15 PD=520e-9 PS=520e-9 NRD=1.16667 NRS=1.16667 M=1
mi13__i19__i4__nm2 n3__i13__i19__i4__net2 n5__i13__net1 n956__vss n640__vss g45n1svt L=45e-9 W=120e-9 AD=16.8e-15 AS=16.8e-15 PD=520e-9 PS=520e-9 NRD=1.16667 NRS=1.16667 M=1
mi13__i19__i4__nm0 n11__i13__net18 i13__i19__i4__net2 n16__i13__net11 n640__vss g45n1svt L=45e-9 W=120e-9 AD=16.8e-15 AS=16.8e-15 PD=520e-9 PS=520e-9 NRD=1.16667 NRS=1.16667 M=1
mi13__i19__i4__nm1 n15__i13__net18 n5__i13__net11 n10__i13__i19__i4__net2 n640__vss g45n1svt L=45e-9 W=120e-9 AD=16.8e-15 AS=16.8e-15 PD=520e-9 PS=520e-9 NRD=1.16667 NRS=1.16667 M=1
mi13__i19__nm0 n8__i13__i19__net1 i13__net1 i13__i19__net3 n640__vss g45n1svt L=45e-9 W=240e-9 AD=33.6e-15 AS=33.6e-15 PD=780e-9 PS=780e-9 NRD=1.16667 NRS=1.16667 M=1
mi13__i19__nm1 i13__i19__net3 i13__net11 n958__vss n640__vss g45n1svt L=45e-9 W=240e-9 AD=38.4e-15 AS=38.4e-15 PD=780e-9 PS=780e-9 NRD=1.16667 NRS=1.16667 M=1
mi13__i19__nm3 n6__i13__net17 i13__i19__net1 n957__vss n640__vss g45n1svt L=45e-9 W=120e-9 AD=16.8e-15 AS=16.8e-15 PD=520e-9 PS=520e-9 NRD=1.16667 NRS=1.16667 M=1
mi13__i17__i4__nm2 n3__i13__i17__i4__net2 n5__i13__a2 n960__vss n640__vss g45n1svt L=45e-9 W=120e-9 AD=16.8e-15 AS=16.8e-15 PD=520e-9 PS=520e-9 NRD=1.16667 NRS=1.16667 M=1
mi13__i17__i4__nm0 n9__i13__net12 i13__i17__i4__net2 n20__i13__a3 n640__vss g45n1svt L=45e-9 W=120e-9 AD=16.8e-15 AS=16.8e-15 PD=520e-9 PS=520e-9 NRD=1.16667 NRS=1.16667 M=1
mi13__i17__i4__nm1 n13__i13__net12 n5__i13__a3 n10__i13__i17__i4__net2 n640__vss g45n1svt L=45e-9 W=120e-9 AD=16.8e-15 AS=16.8e-15 PD=520e-9 PS=520e-9 NRD=1.16667 NRS=1.16667 M=1
mi13__i17__nm0 n8__i13__i17__net1 i13__a2 i13__i17__net3 n640__vss g45n1svt L=45e-9 W=240e-9 AD=33.6e-15 AS=33.6e-15 PD=780e-9 PS=780e-9 NRD=1.16667 NRS=1.16667 M=1
mi13__i17__nm1 i13__i17__net3 i13__a3 n962__vss n640__vss g45n1svt L=45e-9 W=240e-9 AD=38.4e-15 AS=38.4e-15 PD=780e-9 PS=780e-9 NRD=1.16667 NRS=1.16667 M=1
mi13__i17__nm3 n10__i13__net11 i13__i17__net1 n961__vss n640__vss g45n1svt L=45e-9 W=120e-9 AD=16.8e-15 AS=16.8e-15 PD=520e-9 PS=520e-9 NRD=1.16667 NRS=1.16667 M=1
mi13__i18__i4__nm2 n5__i13__i18__i4__net2 n8__i13__net2 n1038__vss n640__vss g45n1svt L=45e-9 W=120e-9 AD=16.8e-15 AS=16.8e-15 PD=520e-9 PS=520e-9 NRD=1.16667 NRS=1.16667 M=1
mi13__i18__i4__nm0 r0 i13__i18__i4__net2 n20__i13__net12 n640__vss g45n1svt L=45e-9 W=120e-9 AD=16.8e-15 AS=16.8e-15 PD=520e-9 PS=520e-9 NRD=1.16667 NRS=1.16667 M=1
mi13__i18__i4__nm1 n8__r0 n8__i13__net12 n8__i13__i18__i4__net2 n640__vss g45n1svt L=45e-9 W=120e-9 AD=16.8e-15 AS=16.8e-15 PD=520e-9 PS=520e-9 NRD=1.16667 NRS=1.16667 M=1
mi13__i18__nm0 n8__i13__i18__net1 n4__i13__net2 i13__i18__net3 n640__vss g45n1svt L=45e-9 W=240e-9 AD=33.6e-15 AS=33.6e-15 PD=780e-9 PS=780e-9 NRD=1.16667 NRS=1.16667 M=1
mi13__i18__nm1 i13__i18__net3 n4__i13__net12 n1040__vss n640__vss g45n1svt L=45e-9 W=240e-9 AD=38.4e-15 AS=38.4e-15 PD=780e-9 PS=780e-9 NRD=1.16667 NRS=1.16667 M=1
mi13__i18__nm3 n10__i13__net7 n4__i13__i18__net1 n1039__vss n640__vss g45n1svt L=45e-9 W=120e-9 AD=16.8e-15 AS=16.8e-15 PD=520e-9 PS=520e-9 NRD=1.16667 NRS=1.16667 M=1
mi13__i16__i4__nm2 n5__i13__i16__i4__net2 n8__i13__a0 n1041__vss n640__vss g45n1svt L=45e-9 W=120e-9 AD=16.8e-15 AS=16.8e-15 PD=520e-9 PS=520e-9 NRD=1.16667 NRS=1.16667 M=1
mi13__i16__i4__nm0 n11__i13__net2 i13__i16__i4__net2 n20__i13__a1 n640__vss g45n1svt L=45e-9 W=120e-9 AD=16.8e-15 AS=16.8e-15 PD=520e-9 PS=520e-9 NRD=1.16667 NRS=1.16667 M=1
mi13__i16__i4__nm1 n18__i13__net2 n8__i13__a1 n8__i13__i16__i4__net2 n640__vss g45n1svt L=45e-9 W=120e-9 AD=16.8e-15 AS=16.8e-15 PD=520e-9 PS=520e-9 NRD=1.16667 NRS=1.16667 M=1
mi13__i16__nm0 n8__i13__i16__net1 n4__i13__a0 i13__i16__net3 n640__vss g45n1svt L=45e-9 W=240e-9 AD=33.6e-15 AS=33.6e-15 PD=780e-9 PS=780e-9 NRD=1.16667 NRS=1.16667 M=1
mi13__i16__nm1 i13__i16__net3 n4__i13__a1 n1043__vss n640__vss g45n1svt L=45e-9 W=240e-9 AD=38.4e-15 AS=38.4e-15 PD=780e-9 PS=780e-9 NRD=1.16667 NRS=1.16667 M=1
mi13__i16__nm3 n12__i13__net1 n4__i13__i16__net1 n1042__vss n640__vss g45n1svt L=45e-9 W=120e-9 AD=16.8e-15 AS=16.8e-15 PD=520e-9 PS=520e-9 NRD=1.16667 NRS=1.16667 M=1
mi13__i15__nm2 n3__i13__i15__net2 n6__x_out_3 n963__vss n640__vss g45n1svt L=45e-9 W=120e-9 AD=16.8e-15 AS=16.8e-15 PD=520e-9 PS=520e-9 NRD=1.16667 NRS=1.16667 M=1
mi13__i15__nm0 n9__i13__a3 i13__i15__net2 n13__y_out_3 n640__vss g45n1svt L=45e-9 W=120e-9 AD=16.8e-15 AS=16.8e-15 PD=520e-9 PS=520e-9 NRD=1.16667 NRS=1.16667 M=1
mi13__i15__nm1 n13__i13__a3 y_out_3 n10__i13__i15__net2 n640__vss g45n1svt L=45e-9 W=120e-9 AD=16.8e-15 AS=16.8e-15 PD=520e-9 PS=520e-9 NRD=1.16667 NRS=1.16667 M=1
mi13__i14__nm2 n3__i13__i14__net2 n6__x_out_2 n964__vss n640__vss g45n1svt L=45e-9 W=120e-9 AD=16.8e-15 AS=16.8e-15 PD=520e-9 PS=520e-9 NRD=1.16667 NRS=1.16667 M=1
mi13__i14__nm0 n9__i13__a2 i13__i14__net2 n12__y_out_2 n640__vss g45n1svt L=45e-9 W=120e-9 AD=16.8e-15 AS=16.8e-15 PD=520e-9 PS=520e-9 NRD=1.16667 NRS=1.16667 M=1
mi13__i14__nm1 n15__i13__a2 y_out_2 n10__i13__i14__net2 n640__vss g45n1svt L=45e-9 W=120e-9 AD=16.8e-15 AS=16.8e-15 PD=520e-9 PS=520e-9 NRD=1.16667 NRS=1.16667 M=1
mi13__i13__nm2 n5__i13__i13__net2 n9__x_out_1 n1058__vss n640__vss g45n1svt L=45e-9 W=120e-9 AD=16.8e-15 AS=16.8e-15 PD=520e-9 PS=520e-9 NRD=1.16667 NRS=1.16667 M=1
mi13__i13__nm0 n9__i13__a1 i13__i13__net2 n12__y_out_1 n640__vss g45n1svt L=45e-9 W=120e-9 AD=16.8e-15 AS=16.8e-15 PD=520e-9 PS=520e-9 NRD=1.16667 NRS=1.16667 M=1
mi13__i13__nm1 n16__i13__a1 n4__y_out_1 n8__i13__i13__net2 n640__vss g45n1svt L=45e-9 W=120e-9 AD=16.8e-15 AS=16.8e-15 PD=520e-9 PS=520e-9 NRD=1.16667 NRS=1.16667 M=1
mi13__i12__nm2 n5__i13__i12__net2 n4__y_out_0 n1059__vss n640__vss g45n1svt L=45e-9 W=120e-9 AD=16.8e-15 AS=16.8e-15 PD=520e-9 PS=520e-9 NRD=1.16667 NRS=1.16667 M=1
mi13__i12__nm0 n9__i13__a0 i13__i12__net2 n14__x_out_0 n640__vss g45n1svt L=45e-9 W=120e-9 AD=16.8e-15 AS=16.8e-15 PD=520e-9 PS=520e-9 NRD=1.16667 NRS=1.16667 M=1
mi13__i12__nm1 n18__i13__a0 n9__x_out_0 n8__i13__i12__net2 n640__vss g45n1svt L=45e-9 W=120e-9 AD=16.8e-15 AS=16.8e-15 PD=520e-9 PS=520e-9 NRD=1.16667 NRS=1.16667 M=1
mi13__nm0 n9__i13__net3 n4__i13__net23 n1037__vss n640__vss g45n1svt L=45e-9 W=120e-9 AD=16.8e-15 AS=16.8e-15 PD=540e-9 PS=540e-9 NRD=1.16667 NRS=1.16667 M=1
mi13__nm1 n1037__vss n4__i13__net17 n4__i13__net3 n640__vss g45n1svt L=45e-9 W=120e-9 AD=19.2e-15 AS=19.2e-15 PD=540e-9 PS=540e-9 NRD=1.16667 NRS=1.16667 M=1
mi13__nm2 n3__r2 n3__i13__net3 n1036__vss n640__vss g45n1svt L=45e-9 W=120e-9 AD=16.8e-15 AS=16.8e-15 PD=520e-9 PS=520e-9 NRD=1.16667 NRS=1.16667 M=1
mi9__i1__nm1_1__rcx n27__shift n5__i9__net1 i9__i1__net1 n640__vss g45n1svt L=45e-9 W=360e-9 AD=57.6e-15 AS=57.6e-15 PD=1.02e-6 PS=1.02e-6 NRD=1.16667 NRS=1.16667 M=1
mi9__i1__nm1 n3__i9__i1__net1 n4__i9__net1 n27__shift n640__vss g45n1svt L=45e-9 W=360e-9 AD=57.6e-15 AS=57.6e-15 PD=1.04e-6 PS=1.04e-6 NRD=1.16667 NRS=1.16667 M=1
mi9__i1__nm0_1__rcx n764__vss n14__ck4 n3__i9__i1__net1 n640__vss g45n1svt L=45e-9 W=360e-9 AD=57.6e-15 AS=57.6e-15 PD=1.04e-6 PS=1.04e-6 NRD=1.16667 NRS=1.16667 M=1
mi9__i1__nm0 n6__i9__i1__net1 n13__ck4 n764__vss n640__vss g45n1svt L=45e-9 W=360e-9 AD=50.4e-15 AS=50.4e-15 PD=1.02e-6 PS=1.02e-6 NRD=1.16667 NRS=1.16667 M=1
mi9__i4__nm0 n12__i9__i4__net1 n2__ck_b n8__ck4 n640__vss g45n1svt L=45e-9 W=120e-9 AD=16.8e-15 AS=16.8e-15 PD=520e-9 PS=520e-9 NRD=1.16667 NRS=1.16667 M=1
mi9__i4__nm8 n805__vss n2__i9__i4__net2 n8__i9__i4__net1 n640__vss g45n1svt L=570e-9 W=120e-9 AD=16.8e-15 AS=16.8e-15 PD=520e-9 PS=520e-9 NRD=1.16667 NRS=1.16667 M=1
mi9__i4__nm18 n804__vss n2__reset_buff n15__i9__i4__net1 n640__vss g45n1svt L=45e-9 W=120e-9 AD=16.8e-15 AS=16.8e-15 PD=520e-9 PS=520e-9 NRD=1.16667 NRS=1.16667 M=1
mi9__i4__nm2_1__rcx n9__i9__i4__net2 n6__i9__i4__net1 n803__vss n640__vss g45n1svt L=45e-9 W=240e-9 AD=38.4e-15 AS=38.4e-15 PD=780e-9 PS=780e-9 NRD=1.16667 NRS=1.16667 M=1
mi9__i4__nm2 n802__vss n5__i9__i4__net1 n9__i9__i4__net2 n640__vss g45n1svt L=45e-9 W=240e-9 AD=33.6e-15 AS=33.6e-15 PD=780e-9 PS=780e-9 NRD=1.16667 NRS=1.16667 M=1
mi9__i4__nm12 n12__i9__i4__net5 n4__ck_buff n10__i9__i4__net2 n640__vss g45n1svt L=45e-9 W=120e-9 AD=16.8e-15 AS=16.8e-15 PD=520e-9 PS=520e-9 NRD=1.16667 NRS=1.16667 M=1
mi9__i4__nm15 n788__vss n2__i9__i4__net4 n8__i9__i4__net5 n640__vss g45n1svt L=570e-9 W=120e-9 AD=16.8e-15 AS=16.8e-15 PD=520e-9 PS=520e-9 NRD=1.16667 NRS=1.16667 M=1
mi9__i4__nm13_1__rcx n8__i9__i4__net4 n6__i9__i4__net5 n783__vss n640__vss g45n1svt L=45e-9 W=240e-9 AD=38.4e-15 AS=38.4e-15 PD=780e-9 PS=780e-9 NRD=1.16667 NRS=1.16667 M=1
mi9__i4__nm13 n778__vss n5__i9__i4__net5 n8__i9__i4__net4 n640__vss g45n1svt L=45e-9 W=240e-9 AD=33.6e-15 AS=33.6e-15 PD=780e-9 PS=780e-9 NRD=1.16667 NRS=1.16667 M=1
mi9__i4__nm16 n6__i9__net2 n6__i9__i4__net4 n777__vss n640__vss g45n1svt L=45e-9 W=240e-9 AD=33.6e-15 AS=33.6e-15 PD=760e-9 PS=760e-9 NRD=1.16667 NRS=1.16667 M=1
mi9__i4__nm17 n9__i9__net1 n4__i9__net2 n772__vss n640__vss g45n1svt L=45e-9 W=240e-9 AD=33.6e-15 AS=33.6e-15 PD=760e-9 PS=760e-9 NRD=1.16667 NRS=1.16667 M=1
mi12__nm2 n11__i12__bcore_bar n11__serial_out n1017__vss n640__vss g45n1svt L=45e-9 W=120e-9 AD=16.8e-15 AS=16.8e-15 PD=520e-9 PS=520e-9 NRD=1.16667 NRS=1.16667 M=1

.ends Top_Level

