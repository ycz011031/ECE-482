** Generated for: hspiceD
** Generated on: Dec  4 22:36:02 2024
** Design library name: ECE482_HW
** Design cell name: Top_Level
** Design view name: schematic


.TEMP 25.0
.OPTION
+    ARTIST=2
+    INGOLD=2
+    PARHIER=LOCAL
+    PSF=2

** Library name: ECE482_HW
** Cell name: inv_1v
** View name: schematic
.subckt inv_1v in out vdd vss
m2 out in vdd vdd g45p1svt L=45e-9 W=240e-9 AD=33.6e-15 AS=33.6e-15 PD=760e-9 PS=760e-9 NRD=583.333e-3 NRS=583.333e-3 M=1
m0 out in vss vss g45n1svt L=45e-9 W=120e-9 AD=16.8e-15 AS=16.8e-15 PD=520e-9 PS=520e-9 NRD=1.16667 NRS=1.16667 M=1
.ends inv_1v
** End of subcircuit definition.

** Library name: ECE482_HW
** Cell name: reg_1b
** View name: schematic
.subckt reg_1b clk clk_b d q q_b rst rstb vdd vss
mnm15 net5 net4 vss vss g45n1svt L=570e-9 W=120e-9 AD=16.8e-15 AS=16.8e-15 PD=520e-9 PS=520e-9 NRD=1.16667 NRS=1.16667 M=1
mnm13 net4 net5 vss vss g45n1svt L=45e-9 W=480e-9 AD=67.2e-15 AS=67.2e-15 PD=1.24e-6 PS=1.24e-6 NRD=291.667e-3 NRS=291.667e-3 M=1
mnm18 net1 rst vss vss g45n1svt L=45e-9 W=120e-9 AD=16.8e-15 AS=16.8e-15 PD=520e-9 PS=520e-9 NRD=1.16667 NRS=1.16667 M=1
mnm8 net1 net2 vss vss g45n1svt L=570e-9 W=120e-9 AD=16.8e-15 AS=16.8e-15 PD=520e-9 PS=520e-9 NRD=1.16667 NRS=1.16667 M=1
mnm16 q_b net4 vss vss g45n1svt L=45e-9 W=240e-9 AD=33.6e-15 AS=33.6e-15 PD=760e-9 PS=760e-9 NRD=583.333e-3 NRS=583.333e-3 M=1
mnm17 q q_b vss vss g45n1svt L=45e-9 W=240e-9 AD=33.6e-15 AS=33.6e-15 PD=760e-9 PS=760e-9 NRD=583.333e-3 NRS=583.333e-3 M=1
mnm2 net2 net1 vss vss g45n1svt L=45e-9 W=480e-9 AD=67.2e-15 AS=67.2e-15 PD=1.24e-6 PS=1.24e-6 NRD=291.667e-3 NRS=291.667e-3 M=1
mnm12 net2 clk net5 vss g45n1svt L=45e-9 W=120e-9 AD=16.8e-15 AS=16.8e-15 PD=520e-9 PS=520e-9 NRD=1.16667 NRS=1.16667 M=1
mnm0 d clk_b net1 vss g45n1svt L=45e-9 W=120e-9 AD=16.8e-15 AS=16.8e-15 PD=520e-9 PS=520e-9 NRD=1.16667 NRS=1.16667 M=1
mpm10 net5 net4 vdd vdd g45p1svt L=180e-9 W=120e-9 AD=16.8e-15 AS=16.8e-15 PD=520e-9 PS=520e-9 NRD=1.16667 NRS=1.16667 M=1
mpm9 net4 net5 vdd vdd g45p1svt L=45e-9 W=960e-9 AD=134.4e-15 AS=134.4e-15 PD=2.2e-6 PS=2.2e-6 NRD=145.833e-3 NRS=145.833e-3 M=1
mpm8 net2 clk_b net5 vdd g45p1svt L=45e-9 W=120e-9 AD=16.8e-15 AS=16.8e-15 PD=520e-9 PS=520e-9 NRD=1.16667 NRS=1.16667 M=1
mpm2 net1 net2 vdd vdd g45p1svt L=180e-9 W=120e-9 AD=16.8e-15 AS=16.8e-15 PD=520e-9 PS=520e-9 NRD=1.16667 NRS=1.16667 M=1
mpm1 net2 net1 vdd vdd g45p1svt L=45e-9 W=960e-9 AD=134.4e-15 AS=134.4e-15 PD=2.2e-6 PS=2.2e-6 NRD=145.833e-3 NRS=145.833e-3 M=1
mpm0 d clk net1 vdd g45p1svt L=45e-9 W=120e-9 AD=16.8e-15 AS=16.8e-15 PD=520e-9 PS=520e-9 NRD=1.16667 NRS=1.16667 M=1
mpm15 net5 rstb vdd vdd g45p1svt L=45e-9 W=120e-9 AD=16.8e-15 AS=16.8e-15 PD=520e-9 PS=520e-9 NRD=1.16667 NRS=1.16667 M=1
mpm13 q q_b vdd vdd g45p1svt L=45e-9 W=480e-9 AD=67.2e-15 AS=67.2e-15 PD=1.24e-6 PS=1.24e-6 NRD=291.667e-3 NRS=291.667e-3 M=1
mpm11 q_b net4 vdd vdd g45p1svt L=45e-9 W=480e-9 AD=67.2e-15 AS=67.2e-15 PD=1.24e-6 PS=1.24e-6 NRD=291.667e-3 NRS=291.667e-3 M=1
.ends reg_1b
** End of subcircuit definition.

** Library name: ECE482_HW
** Cell name: hw10_3_deskew
** View name: schematic
.subckt hw10_3_deskew clk clk_b phi phi_b vdd vss
mnm6 phi_b phi vss vss g45n1svt L=45e-9 W=240e-9 AD=33.6e-15 AS=33.6e-15 PD=760e-9 PS=760e-9 NRD=583.333e-3 NRS=583.333e-3 M=1
mnm5 phi phi_b vss vss g45n1svt L=45e-9 W=240e-9 AD=33.6e-15 AS=33.6e-15 PD=760e-9 PS=760e-9 NRD=583.333e-3 NRS=583.333e-3 M=1
mnm3 phi clk_b vss vss g45n1svt L=45e-9 W=120e-9 AD=16.8e-15 AS=16.8e-15 PD=520e-9 PS=520e-9 NRD=1.16667 NRS=1.16667 M=1
mnm2 vdd clk phi vss g45n1svt L=45e-9 W=120e-9 AD=16.8e-15 AS=16.8e-15 PD=520e-9 PS=520e-9 NRD=1.16667 NRS=1.16667 M=1
mnm1 vdd clk_b phi_b vss g45n1svt L=45e-9 W=120e-9 AD=16.8e-15 AS=16.8e-15 PD=520e-9 PS=520e-9 NRD=1.16667 NRS=1.16667 M=1
mnm0 phi_b clk vss vss g45n1svt L=45e-9 W=120e-9 AD=16.8e-15 AS=16.8e-15 PD=520e-9 PS=520e-9 NRD=1.16667 NRS=1.16667 M=1
mpm6 phi_b phi vdd vdd g45p1svt L=45e-9 W=480e-9 AD=67.2e-15 AS=67.2e-15 PD=1.24e-6 PS=1.24e-6 NRD=291.667e-3 NRS=291.667e-3 M=1
mpm5 phi phi_b vdd vdd g45p1svt L=45e-9 W=480e-9 AD=67.2e-15 AS=67.2e-15 PD=1.24e-6 PS=1.24e-6 NRD=291.667e-3 NRS=291.667e-3 M=1
mpm3 vss clk phi vdd g45p1svt L=45e-9 W=240e-9 AD=33.6e-15 AS=33.6e-15 PD=760e-9 PS=760e-9 NRD=583.333e-3 NRS=583.333e-3 M=1
mpm2 phi clk_b vdd vdd g45p1svt L=45e-9 W=240e-9 AD=33.6e-15 AS=33.6e-15 PD=760e-9 PS=760e-9 NRD=583.333e-3 NRS=583.333e-3 M=1
mpm1 vss clk_b phi_b vdd g45p1svt L=45e-9 W=240e-9 AD=33.6e-15 AS=33.6e-15 PD=760e-9 PS=760e-9 NRD=583.333e-3 NRS=583.333e-3 M=1
mpm0 phi_b clk vdd vdd g45p1svt L=45e-9 W=240e-9 AD=33.6e-15 AS=33.6e-15 PD=760e-9 PS=760e-9 NRD=583.333e-3 NRS=583.333e-3 M=1
.ends hw10_3_deskew
** End of subcircuit definition.

** Library name: ECE482_HW
** Cell name: clk_div4
** View name: schematic
.subckt clk_div4 clk clk_out clk_out_b rst vdd vss
mpm17 clk_out net9 vdd vdd g45p1svt L=45e-9 W=480e-9 AD=67.2e-15 AS=67.2e-15 PD=1.24e-6 PS=1.24e-6 NRD=291.667e-3 NRS=291.667e-3 M=1
mpm1 net6 rst vdd vdd g45p1svt L=45e-9 W=240e-9 AD=33.6e-15 AS=33.6e-15 PD=760e-9 PS=760e-9 NRD=583.333e-3 NRS=583.333e-3 M=1
mpm0 net3 clk vdd vdd g45p1svt L=45e-9 W=240e-9 AD=33.6e-15 AS=33.6e-15 PD=760e-9 PS=760e-9 NRD=583.333e-3 NRS=583.333e-3 M=1
mpm16 clk_out_b net10 vdd vdd g45p1svt L=45e-9 W=480e-9 AD=67.2e-15 AS=67.2e-15 PD=1.24e-6 PS=1.24e-6 NRD=291.667e-3 NRS=291.667e-3 M=1
mnm0 net3 clk vss vss g45n1svt L=45e-9 W=120e-9 AD=16.8e-15 AS=16.8e-15 PD=520e-9 PS=520e-9 NRD=1.16667 NRS=1.16667 M=1
mnm14 clk_out_b net10 vss vss g45n1svt L=45e-9 W=240e-9 AD=33.6e-15 AS=33.6e-15 PD=760e-9 PS=760e-9 NRD=583.333e-3 NRS=583.333e-3 M=1
mnm1 net6 rst vss vss g45n1svt L=45e-9 W=120e-9 AD=16.8e-15 AS=16.8e-15 PD=520e-9 PS=520e-9 NRD=1.16667 NRS=1.16667 M=1
mnm15 clk_out net9 vss vss g45n1svt L=45e-9 W=240e-9 AD=33.6e-15 AS=33.6e-15 PD=760e-9 PS=760e-9 NRD=583.333e-3 NRS=583.333e-3 M=1
xi6 net7 net1 net8 net11 net8 rst net6 vdd vss reg_1b
xi5 clk net3 net1 net7 net1 rst net6 vdd vss reg_1b
xi7 net11 net8 net10 net9 vdd vss hw10_3_deskew
.ends clk_div4
** End of subcircuit definition.

** Library name: ECE482_HW
** Cell name: data_reg_bank
** View name: schematic
.subckt data_reg_bank clk rst vdd vss clk_div4_out clk_div4_out_b x_in_0 x_in_1 x_in_2 x_in_3 x_out_0 x_out_1 x_out_2 x_out_3 x_out_b_0 x_out_b_1 x_out_b_2 x_out_b_3 y_in_0 y_in_1 y_in_2 y_in_3 y_out_0 y_out_1 y_out_2 y_out_3 y_out_b_0 y_out_b_1 y_out_b_2 y_out_b_3
mnm10 clk_div4_out_b net7 vss vss g45n1svt L=45e-9 W=240e-9 AD=33.6e-15 AS=33.6e-15 PD=760e-9 PS=760e-9 NRD=583.333e-3 NRS=583.333e-3 M=1
mnm9 clk_div4_out net11 vss vss g45n1svt L=45e-9 W=240e-9 AD=33.6e-15 AS=33.6e-15 PD=760e-9 PS=760e-9 NRD=583.333e-3 NRS=583.333e-3 M=1
mnm8 net4 rst vss vss g45n1svt L=45e-9 W=1.44e-6 AD=201.6e-15 AS=201.6e-15 PD=3.16e-6 PS=3.16e-6 NRD=97.2222e-3 NRS=97.2222e-3 M=1
mnm7 net3 net4 vss vss g45n1svt L=45e-9 W=1.44e-6 AD=201.6e-15 AS=201.6e-15 PD=3.16e-6 PS=3.16e-6 NRD=97.2222e-3 NRS=97.2222e-3 M=1
mnm1 net10 net11 vss vss g45n1svt L=45e-9 W=1.44e-6 AD=201.6e-15 AS=201.6e-15 PD=3.16e-6 PS=3.16e-6 NRD=97.2222e-3 NRS=97.2222e-3 M=1
mnm0 net9 net7 vss vss g45n1svt L=45e-9 W=1.44e-6 AD=201.6e-15 AS=201.6e-15 PD=3.16e-6 PS=3.16e-6 NRD=97.2222e-3 NRS=97.2222e-3 M=1
mpm10 clk_div4_out_b net7 vdd vdd g45p1svt L=45e-9 W=480e-9 AD=67.2e-15 AS=67.2e-15 PD=1.24e-6 PS=1.24e-6 NRD=291.667e-3 NRS=291.667e-3 M=1
mpm9 clk_div4_out net11 vdd vdd g45p1svt L=45e-9 W=480e-9 AD=67.2e-15 AS=67.2e-15 PD=1.24e-6 PS=1.24e-6 NRD=291.667e-3 NRS=291.667e-3 M=1
mpm8 net4 rst vdd vdd g45p1svt L=45e-9 W=2.88e-6 AD=403.2e-15 AS=403.2e-15 PD=6.04e-6 PS=6.04e-6 NRD=48.6111e-3 NRS=48.6111e-3 M=1
mpm7 net3 net4 vdd vdd g45p1svt L=45e-9 W=2.88e-6 AD=403.2e-15 AS=403.2e-15 PD=6.04e-6 PS=6.04e-6 NRD=48.6111e-3 NRS=48.6111e-3 M=1
mpm3 net10 net11 vdd vdd g45p1svt L=45e-9 W=2.88e-6 AD=403.2e-15 AS=403.2e-15 PD=6.04e-6 PS=6.04e-6 NRD=48.6111e-3 NRS=48.6111e-3 M=1
mpm2 net9 net7 vdd vdd g45p1svt L=45e-9 W=2.88e-6 AD=403.2e-15 AS=403.2e-15 PD=6.04e-6 PS=6.04e-6 NRD=48.6111e-3 NRS=48.6111e-3 M=1
xi16 net10 net9 y_in_0 y_out_0 y_out_b_0 net3 net4 vdd vss reg_1b
xi15 net10 net9 y_in_1 y_out_1 y_out_b_1 net3 net4 vdd vss reg_1b
xi14 net10 net9 y_in_2 y_out_2 y_out_b_2 net3 net4 vdd vss reg_1b
xi13 net10 net9 y_in_3 y_out_3 y_out_b_3 net3 net4 vdd vss reg_1b
xi12 net10 net9 x_in_0 x_out_0 x_out_b_0 net3 net4 vdd vss reg_1b
xi11 net10 net9 x_in_1 x_out_1 x_out_b_1 net3 net4 vdd vss reg_1b
xi10 net10 net9 x_in_2 x_out_2 x_out_b_2 net3 net4 vdd vss reg_1b
xi9 net10 net9 x_in_3 x_out_3 x_out_b_3 net3 net4 vdd vss reg_1b
xi17 clk net7 net11 rst vdd vss clk_div4
.ends data_reg_bank
** End of subcircuit definition.

** Library name: ECE482_HW
** Cell name: intergrated
** View name: schematic
.subckt intergrated a b clk clk_b q q_b rst rstb shift vdd vss
mnm21 net79 shift vss vss g45n1svt L=45e-9 W=120e-9 AD=16.8e-15 AS=16.8e-15 PD=520e-9 PS=520e-9 NRD=1.16667 NRS=1.16667 M=1
mnm20 b net79 net73 vss g45n1svt L=45e-9 W=120e-9 AD=16.8e-15 AS=16.8e-15 PD=520e-9 PS=520e-9 NRD=1.16667 NRS=1.16667 M=1
mnm22 a shift net73 vss g45n1svt L=45e-9 W=120e-9 AD=16.8e-15 AS=16.8e-15 PD=520e-9 PS=520e-9 NRD=1.16667 NRS=1.16667 M=1
mnm12 net75 clk net76 vss g45n1svt L=45e-9 W=120e-9 AD=16.8e-15 AS=16.8e-15 PD=520e-9 PS=520e-9 NRD=1.16667 NRS=1.16667 M=1
mnm0 net73 clk_b net74 vss g45n1svt L=45e-9 W=120e-9 AD=16.8e-15 AS=16.8e-15 PD=520e-9 PS=520e-9 NRD=1.16667 NRS=1.16667 M=1
mnm13 net77 net76 vss vss g45n1svt L=45e-9 W=480e-9 AD=67.2e-15 AS=67.2e-15 PD=1.24e-6 PS=1.24e-6 NRD=291.667e-3 NRS=291.667e-3 M=1
mnm16 q_b net77 vss vss g45n1svt L=45e-9 W=240e-9 AD=33.6e-15 AS=33.6e-15 PD=760e-9 PS=760e-9 NRD=583.333e-3 NRS=583.333e-3 M=1
mnm2 net75 net74 vss vss g45n1svt L=45e-9 W=480e-9 AD=67.2e-15 AS=67.2e-15 PD=1.24e-6 PS=1.24e-6 NRD=291.667e-3 NRS=291.667e-3 M=1
mnm17 q q_b vss vss g45n1svt L=45e-9 W=240e-9 AD=33.6e-15 AS=33.6e-15 PD=760e-9 PS=760e-9 NRD=583.333e-3 NRS=583.333e-3 M=1
mnm15 net76 net77 vss vss g45n1svt L=570e-9 W=120e-9 AD=16.8e-15 AS=16.8e-15 PD=520e-9 PS=520e-9 NRD=1.16667 NRS=1.16667 M=1
mnm18 net74 rst vss vss g45n1svt L=45e-9 W=120e-9 AD=16.8e-15 AS=16.8e-15 PD=520e-9 PS=520e-9 NRD=1.16667 NRS=1.16667 M=1
mnm8 net74 net75 vss vss g45n1svt L=570e-9 W=120e-9 AD=16.8e-15 AS=16.8e-15 PD=520e-9 PS=520e-9 NRD=1.16667 NRS=1.16667 M=1
mpm18 net79 shift vdd vdd g45p1svt L=45e-9 W=240e-9 AD=33.6e-15 AS=33.6e-15 PD=760e-9 PS=760e-9 NRD=583.333e-3 NRS=583.333e-3 M=1
mpm19 b shift net73 vdd g45p1svt L=45e-9 W=240e-9 AD=33.6e-15 AS=33.6e-15 PD=760e-9 PS=760e-9 NRD=583.333e-3 NRS=583.333e-3 M=1
mpm16 a net79 net73 vdd g45p1svt L=45e-9 W=240e-9 AD=33.6e-15 AS=33.6e-15 PD=760e-9 PS=760e-9 NRD=583.333e-3 NRS=583.333e-3 M=1
mpm8 net75 clk_b net76 vdd g45p1svt L=45e-9 W=120e-9 AD=16.8e-15 AS=16.8e-15 PD=520e-9 PS=520e-9 NRD=1.16667 NRS=1.16667 M=1
mpm0 net73 clk net74 vdd g45p1svt L=45e-9 W=120e-9 AD=16.8e-15 AS=16.8e-15 PD=520e-9 PS=520e-9 NRD=1.16667 NRS=1.16667 M=1
mpm15 net76 rstb vdd vdd g45p1svt L=45e-9 W=120e-9 AD=16.8e-15 AS=16.8e-15 PD=520e-9 PS=520e-9 NRD=1.16667 NRS=1.16667 M=1
mpm9 net77 net76 vdd vdd g45p1svt L=45e-9 W=960e-9 AD=134.4e-15 AS=134.4e-15 PD=2.2e-6 PS=2.2e-6 NRD=145.833e-3 NRS=145.833e-3 M=1
mpm1 net75 net74 vdd vdd g45p1svt L=45e-9 W=960e-9 AD=134.4e-15 AS=134.4e-15 PD=2.2e-6 PS=2.2e-6 NRD=145.833e-3 NRS=145.833e-3 M=1
mpm11 q_b net77 vdd vdd g45p1svt L=45e-9 W=480e-9 AD=67.2e-15 AS=67.2e-15 PD=1.24e-6 PS=1.24e-6 NRD=291.667e-3 NRS=291.667e-3 M=1
mpm13 q q_b vdd vdd g45p1svt L=45e-9 W=480e-9 AD=67.2e-15 AS=67.2e-15 PD=1.24e-6 PS=1.24e-6 NRD=291.667e-3 NRS=291.667e-3 M=1
mpm10 net76 net77 vdd vdd g45p1svt L=180e-9 W=120e-9 AD=16.8e-15 AS=16.8e-15 PD=520e-9 PS=520e-9 NRD=1.16667 NRS=1.16667 M=1
mpm2 net74 net75 vdd vdd g45p1svt L=180e-9 W=120e-9 AD=16.8e-15 AS=16.8e-15 PD=520e-9 PS=520e-9 NRD=1.16667 NRS=1.16667 M=1
.ends intergrated
** End of subcircuit definition.

** Library name: ECE482_HW
** Cell name: PISO
** View name: schematic
.subckt PISO clk clk_b rst rstb shift serial_out vdd vss r0 r1 r2
xi2 net2 r0 clk clk_b serial_out net5 rst rstb shift vdd vss intergrated
xi1 net1 r1 clk clk_b net2 net4 rst rstb shift vdd vss intergrated
xi0 vss r2 clk clk_b net1 net3 rst rstb shift vdd vss intergrated
.ends PISO
** End of subcircuit definition.

** Library name: ECE482_HW
** Cell name: NAND
** View name: schematic
.subckt NAND a b out vdd vss
mnm1 net1 b vss vss g45n1svt L=45e-9 W=120e-9 AD=16.8e-15 AS=16.8e-15 PD=520e-9 PS=520e-9 NRD=1.16667 NRS=1.16667 M=1
mnm0 out a net1 vss g45n1svt L=45e-9 W=120e-9 AD=16.8e-15 AS=16.8e-15 PD=520e-9 PS=520e-9 NRD=1.16667 NRS=1.16667 M=1
mpm1 out b vdd vdd g45p1svt L=45e-9 W=240e-9 AD=33.6e-15 AS=33.6e-15 PD=760e-9 PS=760e-9 NRD=583.333e-3 NRS=583.333e-3 M=1
mpm0 out a vdd vdd g45p1svt L=45e-9 W=240e-9 AD=33.6e-15 AS=33.6e-15 PD=760e-9 PS=760e-9 NRD=583.333e-3 NRS=583.333e-3 M=1
.ends NAND
** End of subcircuit definition.

** Library name: ECE482_HW
** Cell name: Shift_Signal
** View name: schematic
.subckt Shift_Signal clk clk_b clk_out rst rstb shift vdd vss
xi4 clk clk_b clk_out net1 net2 rst rstb vdd vss reg_1b
xi1 net1 clk_out shift vdd vss NAND
.ends Shift_Signal
** End of subcircuit definition.

** Library name: ECE482_HW
** Cell name: Off_chip_Driver
** View name: schematic
.subckt Off_chip_Driver in out vdd vss
m15 out net5 vss vss g45n2svt L=150e-9 W=600e-6 AD=60e-12 AS=61e-12 PD=612e-6 PS=632.2e-6 NRD=166.667e-6 NRS=169.444e-6 M=1
m14 net5 net4 vss vss g45n2svt L=150e-9 W=166.6e-6 AD=17.15e-12 AS=17.15e-12 PD=179.9e-6 PS=179.9e-6 NRD=617.894e-6 NRS=617.894e-6 M=1
m3 net4 net3 vss vss g45n2svt L=150e-9 W=45.85e-6 AD=5.0435e-12 AS=5.0435e-12 PD=56.12e-6 PS=56.12e-6 NRD=2.39913e-3 NRS=2.39913e-3 M=1
m2 net3 net2 vss vss g45n2svt L=150e-9 W=12.64e-6 AD=1.264e-12 AS=1.896e-12 PD=13.04e-6 PS=25.88e-6 NRD=7.91139e-3 NRS=11.8671e-3 M=1
m1 net2 net1 vss vss g45n2svt L=150e-9 W=3.48e-6 AD=522e-15 AS=522e-15 PD=7.26e-6 PS=7.26e-6 NRD=43.1034e-3 NRS=43.1034e-3 M=1
m0 net1 in vss vss g45n2svt L=150e-9 W=960e-9 AD=144e-15 AS=144e-15 PD=2.22e-6 PS=2.22e-6 NRD=156.25e-3 NRS=156.25e-3 M=1
m17 out net5 vdd vdd g45p2svt L=150e-9 W=822e-6 AD=82.2e-12 AS=83.022e-12 PD=842e-6 PS=858.64e-6 NRD=121.655e-6 NRS=122.871e-6 M=1
m16 net5 net4 vdd vdd g45p2svt L=150e-9 W=229.54e-6 AD=23.453e-12 AS=23.453e-12 PD=244.22e-6 PS=244.22e-6 NRD=445.125e-6 NRS=445.125e-6 M=1
m9 net4 net3 vdd vdd g45p2svt L=150e-9 W=62.8e-6 AD=6.28e-12 AS=6.908e-12 PD=64.8e-6 PS=77.56e-6 NRD=1.59236e-3 NRS=1.75159e-3 M=1
m8 net3 net2 vdd vdd g45p2svt L=150e-9 W=17.32e-6 AD=1.732e-12 AS=2.165e-12 PD=18.12e-6 PS=26.98e-6 NRD=5.77367e-3 NRS=7.21709e-3 M=1
m7 net2 net1 vdd vdd g45p2svt L=150e-9 W=4.76e-6 AD=714e-15 AS=714e-15 PD=9.82e-6 PS=9.82e-6 NRD=31.5126e-3 NRS=31.5126e-3 M=1
m6 net1 in vdd vdd g45p2svt L=150e-9 W=1.32e-6 AD=198e-15 AS=198e-15 PD=2.94e-6 PS=2.94e-6 NRD=113.636e-3 NRS=113.636e-3 M=1
.ends Off_chip_Driver
** End of subcircuit definition.

** Library name: ECE482_HW
** Cell name: Level_Shifter_Project
** View name: schematic
.subckt Level_Shifter_Project bio bio_bar bcore vdd vddio vss
mpm0 bcore_bar bcore vdd vdd g45p1svt L=45e-9 W=240e-9 AD=33.6e-15 AS=33.6e-15 PD=760e-9 PS=760e-9 NRD=583.333e-3 NRS=583.333e-3 M=1
m1 bio_bar bio vddio vddio g45p2svt L=150e-9 W=320e-9 AD=48e-15 AS=48e-15 PD=940e-9 PS=940e-9 NRD=468.75e-3 NRS=468.75e-3 M=1
m0 bio bio_bar vddio vddio g45p2svt L=150e-9 W=320e-9 AD=48e-15 AS=48e-15 PD=940e-9 PS=940e-9 NRD=468.75e-3 NRS=468.75e-3 M=1
mnm1 bio_bar bcore vss vss g45n2svt L=150e-9 W=320e-9 AD=48e-15 AS=48e-15 PD=940e-9 PS=940e-9 NRD=468.75e-3 NRS=468.75e-3 M=1
mnm0 bio bcore_bar vss vss g45n2svt L=150e-9 W=320e-9 AD=48e-15 AS=48e-15 PD=940e-9 PS=940e-9 NRD=468.75e-3 NRS=468.75e-3 M=1
mnm2 bcore_bar bcore vss vss g45n1svt L=45e-9 W=120e-9 AD=16.8e-15 AS=16.8e-15 PD=520e-9 PS=520e-9 NRD=1.16667 NRS=1.16667 M=1
.ends Level_Shifter_Project
** End of subcircuit definition.

** Library name: ECE482_HW
** Cell name: xor_tran
** View name: schematic
.subckt xor_tran a b out vdd vss
mpm2 net2 a vdd vdd g45p1svt L=45e-9 W=120e-9 AD=16.8e-15 AS=16.8e-15 PD=520e-9 PS=520e-9 NRD=1.16667 NRS=1.16667 M=1
mpm1 out b a vdd g45p1svt L=45e-9 W=120e-9 AD=16.8e-15 AS=16.8e-15 PD=520e-9 PS=520e-9 NRD=1.16667 NRS=1.16667 M=1
mpm0 b a out vdd g45p1svt L=45e-9 W=120e-9 AD=16.8e-15 AS=16.8e-15 PD=520e-9 PS=520e-9 NRD=1.16667 NRS=1.16667 M=1
mnm2 net2 a vss vss g45n1svt L=45e-9 W=120e-9 AD=16.8e-15 AS=16.8e-15 PD=520e-9 PS=520e-9 NRD=1.16667 NRS=1.16667 M=1
mnm1 out b net2 vss g45n1svt L=45e-9 W=120e-9 AD=16.8e-15 AS=16.8e-15 PD=520e-9 PS=520e-9 NRD=1.16667 NRS=1.16667 M=1
mnm0 b net2 out vss g45n1svt L=45e-9 W=120e-9 AD=16.8e-15 AS=16.8e-15 PD=520e-9 PS=520e-9 NRD=1.16667 NRS=1.16667 M=1
.ends xor_tran
** End of subcircuit definition.

** Library name: ECE482_HW
** Cell name: half_adder
** View name: schematic
.subckt half_adder a b cout sum vdd vss
mpm2 cout net1 vdd vdd g45p1svt L=45e-9 W=120e-9 AD=16.8e-15 AS=16.8e-15 PD=520e-9 PS=520e-9 NRD=1.16667 NRS=1.16667 M=1
mpm0 net1 a vdd vdd g45p1svt L=45e-9 W=120e-9 AD=16.8e-15 AS=16.8e-15 PD=520e-9 PS=520e-9 NRD=1.16667 NRS=1.16667 M=1
mpm1 net1 b vdd vdd g45p1svt L=45e-9 W=120e-9 AD=16.8e-15 AS=16.8e-15 PD=520e-9 PS=520e-9 NRD=1.16667 NRS=1.16667 M=1
mnm3 cout net1 vss vss g45n1svt L=45e-9 W=120e-9 AD=16.8e-15 AS=16.8e-15 PD=520e-9 PS=520e-9 NRD=1.16667 NRS=1.16667 M=1
mnm1 net3 b vss vss g45n1svt L=45e-9 W=120e-9 AD=16.8e-15 AS=16.8e-15 PD=520e-9 PS=520e-9 NRD=1.16667 NRS=1.16667 M=1
mnm0 net1 a net3 vss g45n1svt L=45e-9 W=120e-9 AD=16.8e-15 AS=16.8e-15 PD=520e-9 PS=520e-9 NRD=1.16667 NRS=1.16667 M=1
xi4 a b sum vdd vss xor_tran
.ends half_adder
** End of subcircuit definition.

** Library name: ECE482_HW
** Cell name: adder_circuit
** View name: schematic
.subckt adder_circuit vdd vss r0 r1 r2 x0 x1 x2 x3 y0 y1 y2 y3
mpm2 r2 net3 vdd vdd g45p1svt L=45e-9 W=120e-9 AD=16.8e-15 AS=16.8e-15 PD=520e-9 PS=520e-9 NRD=1.16667 NRS=1.16667 M=1
mpm1 net3 net17 net6 vdd g45p1svt L=45e-9 W=120e-9 AD=16.8e-15 AS=16.8e-15 PD=520e-9 PS=520e-9 NRD=1.16667 NRS=1.16667 M=1
mpm0 net6 net23 vdd vdd g45p1svt L=45e-9 W=120e-9 AD=16.8e-15 AS=16.8e-15 PD=520e-9 PS=520e-9 NRD=1.16667 NRS=1.16667 M=1
mnm2 r2 net3 vss vss g45n1svt L=45e-9 W=120e-9 AD=16.8e-15 AS=16.8e-15 PD=520e-9 PS=520e-9 NRD=1.16667 NRS=1.16667 M=1
mnm1 net3 net17 vss vss g45n1svt L=45e-9 W=120e-9 AD=16.8e-15 AS=16.8e-15 PD=520e-9 PS=520e-9 NRD=1.16667 NRS=1.16667 M=1
mnm0 net3 net23 vss vss g45n1svt L=45e-9 W=120e-9 AD=16.8e-15 AS=16.8e-15 PD=520e-9 PS=520e-9 NRD=1.16667 NRS=1.16667 M=1
xi15 x3 y3 a3 vdd vss xor_tran
xi14 x2 y2 a2 vdd vss xor_tran
xi13 x1 y1 a1 vdd vss xor_tran
xi12 x0 y0 a0 vdd vss xor_tran
xi20 net18 net7 net23 r1 vdd vss half_adder
xi19 net1 net11 net17 net18 vdd vss half_adder
xi18 net2 net12 net7 r0 vdd vss half_adder
xi17 a2 a3 net11 net12 vdd vss half_adder
xi16 a0 a1 net1 net2 vdd vss half_adder
.ends adder_circuit
** End of subcircuit definition.

** Library name: ECE482_HW
** Cell name: Top_Level
** View name: schematic
xi17 reset reset_b vdd vss inv_1v
xi16 ck ck_b vdd vss inv_1v
xi14 ck reset vdd vss ck4 ck4_b x0 x1 x2 x3 x_out_0 x_out_1 x_out_2 x_out_3 x_out_b_0 x_out_b_1 x_out_b_2 x_out_b_3 y0 y1 y2 y3 y_out_0 y_out_1 y_out_2 y_out_3 y_out_b_0 y_out_b_1 y_out_b_2 y_out_b_3 data_reg_bank
xi8 ck ck_b reset reset_b shift serial_out vdd vss r0 r1 r2 PISO
xi9 ck ck_b ck4 reset reset_b shift vdd vss Shift_Signal
xi18 serial_out_high r_out vddio vss Off_chip_Driver
xi12 serial_out_high serial_out_b_high serial_out vdd vddio vss Level_Shifter_Project
xi13 vdd vss r0 r1 r2 x_out_0 x_out_1 x_out_2 x_out_3 y_out_0 y_out_1 y_out_2 y_out_3 adder_circuit
.END
